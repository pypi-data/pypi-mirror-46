(lp0
(ccopy_reg
_reconstructor
p1
(cpygments.token
_TokenType
p2
c__builtin__
tuple
p3
(S'Keyword'
p4
tp5
tp6
Rp7
(dp8
S'parent'
p9
g1
(g2
g3
(ttp10
Rp11
(dp12
S'Number'
p13
g1
(g2
g3
(S'Literal'
p14
g13
tp15
tp16
Rp17
(dp18
S'Integer'
p19
g1
(g2
g3
(g14
g13
g19
tp20
tp21
Rp22
(dp23
g9
g17
sS'Long'
p24
g1
(g2
g3
(g14
g13
g19
g24
tp25
tp26
Rp27
(dp28
g9
g22
sS'subtypes'
p29
c__builtin__
set
p30
((lp31
tp32
Rp33
sbsg29
g30
((lp34
g27
atp35
Rp36
sbsg9
g1
(g2
g3
(g14
tp37
tp38
Rp39
(dp40
S'Scalar'
p41
g1
(g2
g3
(g14
g41
tp42
tp43
Rp44
(dp45
g9
g39
sg29
g30
((lp46
g1
(g2
g3
(g14
g41
S'Plain'
p47
tp48
tp49
Rp50
(dp51
g9
g44
sg29
g30
((lp52
tp53
Rp54
sbatp55
Rp56
sg47
g50
sbsg13
g17
sg9
g11
sS'Other'
p57
g1
(g2
g3
(g14
g57
tp58
tp59
Rp60
(dp61
g9
g39
sg29
g30
((lp62
tp63
Rp64
sbsS'Char'
p65
g1
(g2
g3
(g14
g65
tp66
tp67
Rp68
(dp69
g9
g39
sg29
g30
((lp70
tp71
Rp72
sbsS'String'
p73
g1
(g2
g3
(g14
g73
tp74
tp75
Rp76
(dp77
g65
g1
(g2
g3
(g14
g73
g65
tp78
tp79
Rp80
(dp81
g9
g76
sg29
g30
((lp82
tp83
Rp84
sbsS'Backtick'
p85
g1
(g2
g3
(g14
g73
g85
tp86
tp87
Rp88
(dp89
g9
g76
sg29
g30
((lp90
tp91
Rp92
sbsS'Heredoc'
p93
g1
(g2
g3
(g14
g73
g93
tp94
tp95
Rp96
(dp97
g9
g76
sg29
g30
((lp98
tp99
Rp100
sbsS'Symbol'
p101
g1
(g2
g3
(g14
g73
g101
tp102
tp103
Rp104
(dp105
g9
g76
sg29
g30
((lp106
tp107
Rp108
sbsS'Interpol'
p109
g1
(g2
g3
(g14
g73
g109
tp110
tp111
Rp112
(dp113
g9
g76
sg29
g30
((lp114
tp115
Rp116
sbsS'Delimiter'
p117
g1
(g2
g3
(g14
g73
g117
tp118
tp119
Rp120
(dp121
g9
g76
sg29
g30
((lp122
tp123
Rp124
sbsS'Boolean'
p125
g1
(g2
g3
(g14
g73
g125
tp126
tp127
Rp128
(dp129
g9
g76
sg29
g30
((lp130
tp131
Rp132
sbsS'Character'
p133
g1
(g2
g3
(g14
g73
g133
tp134
tp135
Rp136
(dp137
g9
g76
sg29
g30
((lp138
tp139
Rp140
sbsS'Double'
p141
g1
(g2
g3
(g14
g73
g141
tp142
tp143
Rp144
(dp145
g9
g76
sg29
g30
((lp146
tp147
Rp148
sbsS'Delimeter'
p149
g1
(g2
g3
(g14
g73
g149
tp150
tp151
Rp152
(dp153
g9
g76
sg29
g30
((lp154
tp155
Rp156
sbsS'Atom'
p157
g1
(g2
g3
(g14
g73
g157
tp158
tp159
Rp160
(dp161
g9
g76
sg29
g30
((lp162
tp163
Rp164
sbsS'Affix'
p165
g1
(g2
g3
(g14
g73
g165
tp166
tp167
Rp168
(dp169
g9
g76
sg29
g30
((lp170
tp171
Rp172
sbsS'Name'
p173
g1
(g2
g3
(g14
g73
g173
tp174
tp175
Rp176
(dp177
g9
g76
sg29
g30
((lp178
tp179
Rp180
sbsS'Regex'
p181
g1
(g2
g3
(g14
g73
g181
tp182
tp183
Rp184
(dp185
g9
g76
sg29
g30
((lp186
tp187
Rp188
sbsS'Interp'
p189
g1
(g2
g3
(g14
g73
g189
tp190
tp191
Rp192
(dp193
g9
g76
sg29
g30
((lp194
tp195
Rp196
sbsS'Escape'
p197
g1
(g2
g3
(g14
g73
g197
tp198
tp199
Rp200
(dp201
g9
g76
sg29
g30
((lp202
tp203
Rp204
sbsg29
g30
((lp205
g120
ag104
ag184
ag1
(g2
g3
(g14
g73
S'Doc'
p206
tp207
tp208
Rp209
(dp210
g9
g76
sg29
g30
((lp211
tp212
Rp213
sbag136
ag128
ag144
ag112
ag160
ag152
ag176
ag200
ag1
(g2
g3
(g14
g73
S'Single'
p214
tp215
tp216
Rp217
(dp218
g9
g76
sg29
g30
((lp219
tp220
Rp221
sbag1
(g2
g3
(g14
g73
g57
tp222
tp223
Rp224
(dp225
g9
g76
sg29
g30
((lp226
tp227
Rp228
sbag192
ag88
ag168
ag1
(g2
g3
(g14
g73
S'Moment'
p229
tp230
tp231
Rp232
(dp233
g9
g76
sg29
g30
((lp234
tp235
Rp236
sbag80
ag96
atp237
Rp238
sg214
g217
sg229
g232
sg9
g39
sg57
g224
sg206
g209
sbsg29
g30
((lp239
g76
ag68
ag60
ag1
(g2
g3
(g14
S'Date'
p240
tp241
tp242
Rp243
(dp244
g9
g39
sg29
g30
((lp245
tp246
Rp247
sbag44
ag17
atp248
Rp249
sg240
g243
sbsS'Bin'
p250
g1
(g2
g3
(g14
g13
g250
tp251
tp252
Rp253
(dp254
g9
g17
sg29
g30
((lp255
tp256
Rp257
sbsS'Radix'
p258
g1
(g2
g3
(g14
g13
g258
tp259
tp260
Rp261
(dp262
g9
g17
sg29
g30
((lp263
tp264
Rp265
sbsS'Oct'
p266
g1
(g2
g3
(g14
g13
g266
tp267
tp268
Rp269
(dp270
g9
g17
sg29
g30
((lp271
tp272
Rp273
sbsS'Dec'
p274
g1
(g2
g3
(g14
g13
g274
tp275
tp276
Rp277
(dp278
g9
g17
sg29
g30
((lp279
tp280
Rp281
sbsS'Hex'
p282
g1
(g2
g3
(g14
g13
g282
tp283
tp284
Rp285
(dp286
g9
g17
sg29
g30
((lp287
tp288
Rp289
sbsg29
g30
((lp290
g22
ag261
ag277
ag1
(g2
g3
(g14
g13
S'Decimal'
p291
tp292
tp293
Rp294
(dp295
g9
g17
sg29
g30
((lp296
tp297
Rp298
sbag253
ag1
(g2
g3
(g14
g13
S'Float'
p299
tp300
tp301
Rp302
(dp303
g9
g17
sg29
g30
((lp304
tp305
Rp306
sbag269
ag285
atp307
Rp308
sg291
g294
sg299
g302
sbsS'Generic'
p309
g1
(g2
g3
(g309
tp310
tp311
Rp312
(dp313
g9
g11
sS'Deleted'
p314
g1
(g2
g3
(g309
g314
tp315
tp316
Rp317
(dp318
g9
g312
sg29
g30
((lp319
tp320
Rp321
sbsS'Subheading'
p322
g1
(g2
g3
(g309
g322
tp323
tp324
Rp325
(dp326
g9
g312
sg29
g30
((lp327
tp328
Rp329
sbsS'Heading'
p330
g1
(g2
g3
(g309
g330
tp331
tp332
Rp333
(dp334
g9
g312
sg29
g30
((lp335
tp336
Rp337
sbsS'Emph'
p338
g1
(g2
g3
(g309
g338
tp339
tp340
Rp341
(dp342
g9
g312
sg29
g30
((lp343
tp344
Rp345
sbsS'Prompt'
p346
g1
(g2
g3
(g309
g346
tp347
tp348
Rp349
(dp350
g9
g312
sg29
g30
((lp351
tp352
Rp353
sbsS'Inserted'
p354
g1
(g2
g3
(g309
g354
tp355
tp356
Rp357
(dp358
g9
g312
sg29
g30
((lp359
tp360
Rp361
sbsS'Strong'
p362
g1
(g2
g3
(g309
g362
tp363
tp364
Rp365
(dp366
g9
g312
sg29
g30
((lp367
tp368
Rp369
sbsS'Error'
p370
g1
(g2
g3
(g309
g370
tp371
tp372
Rp373
(dp374
g9
g312
sg29
g30
((lp375
tp376
Rp377
sbsS'Traceback'
p378
g1
(g2
g3
(g309
g378
tp379
tp380
Rp381
(dp382
g9
g312
sg29
g30
((lp383
tp384
Rp385
sbsg29
g30
((lp386
g333
ag325
ag1
(g2
g3
(g309
S'Output'
p387
tp388
tp389
Rp390
(dp391
g9
g312
sg29
g30
((lp392
tp393
Rp394
sbag365
ag341
ag373
ag381
ag357
ag349
ag317
atp395
Rp396
sg387
g390
sbsS'Operator'
p397
g1
(g2
g3
(g397
tp398
tp399
Rp400
(dp401
g9
g11
sS'DBS'
p402
g1
(g2
g3
(g397
g402
tp403
tp404
Rp405
(dp406
g9
g400
sg29
g30
((lp407
tp408
Rp409
sbsg29
g30
((lp410
g405
ag1
(g2
g3
(g397
S'Word'
p411
tp412
tp413
Rp414
(dp415
g9
g400
sg29
g30
((lp416
tp417
Rp418
sbatp419
Rp420
sg411
g414
sbsg73
g76
sg173
g1
(g2
g3
(g173
tp421
tp422
Rp423
(dp424
S'Variable'
p425
g1
(g2
g3
(g173
g425
tp426
tp427
Rp428
(dp429
g9
g423
sS'Class'
p430
g1
(g2
g3
(g173
g425
g430
tp431
tp432
Rp433
(dp434
g9
g428
sg29
g30
((lp435
tp436
Rp437
sbsS'Anonymous'
p438
g1
(g2
g3
(g173
g425
g438
tp439
tp440
Rp441
(dp442
g9
g428
sg29
g30
((lp443
tp444
Rp445
sbsS'Instance'
p446
g1
(g2
g3
(g173
g425
g446
tp447
tp448
Rp449
(dp450
g9
g428
sg29
g30
((lp451
tp452
Rp453
sbsS'Global'
p454
g1
(g2
g3
(g173
g425
g454
tp455
tp456
Rp457
(dp458
g9
g428
sg29
g30
((lp459
tp460
Rp461
sbsg29
g30
((lp462
g441
ag449
ag1
(g2
g3
(g173
g425
S'Magic'
p463
tp464
tp465
Rp466
(dp467
g9
g428
sg29
g30
((lp468
tp469
Rp470
sbag457
ag433
atp471
Rp472
sg463
g466
sbsg397
g1
(g2
g3
(g173
g397
tp473
tp474
Rp475
(dp476
g9
g423
sg29
g30
((lp477
tp478
Rp479
sbsS'Decorator'
p480
g1
(g2
g3
(g173
g480
tp481
tp482
Rp483
(dp484
g9
g423
sg29
g30
((lp485
tp486
Rp487
sbsS'Entity'
p488
g1
(g2
g3
(g173
g488
tp489
tp490
Rp491
(dp492
g9
g423
sg402
g1
(g2
g3
(g173
g488
g402
tp493
tp494
Rp495
(dp496
g9
g491
sg29
g30
((lp497
tp498
Rp499
sbsg29
g30
((lp500
g495
atp501
Rp502
sbsg101
g1
(g2
g3
(g173
g101
tp503
tp504
Rp505
(dp506
g9
g423
sg29
g30
((lp507
tp508
Rp509
sbsS'Property'
p510
g1
(g2
g3
(g173
g510
tp511
tp512
Rp513
(dp514
g9
g423
sg29
g30
((lp515
tp516
Rp517
sbsS'Pseudo'
p518
g1
(g2
g3
(g173
g518
tp519
tp520
Rp521
(dp522
g9
g423
sg29
g30
((lp523
tp524
Rp525
sbsS'Type'
p526
g1
(g2
g3
(g173
g526
tp527
tp528
Rp529
(dp530
g9
g423
sg29
g30
((lp531
tp532
Rp533
sbsS'Classes'
p534
g1
(g2
g3
(g173
g534
tp535
tp536
Rp537
(dp538
g9
g423
sg29
g30
((lp539
tp540
Rp541
sbsS'Tag'
p542
g1
(g2
g3
(g173
g542
tp543
tp544
Rp545
(dp546
g9
g423
sg29
g30
((lp547
tp548
Rp549
sbsS'Constant'
p550
g1
(g2
g3
(g173
g550
tp551
tp552
Rp553
(dp554
g9
g423
sg29
g30
((lp555
tp556
Rp557
sbsS'Function'
p558
g1
(g2
g3
(g173
g558
tp559
tp560
Rp561
(dp562
g9
g423
sg29
g30
((lp563
g1
(g2
g3
(g173
g558
g463
tp564
tp565
Rp566
(dp567
g9
g561
sg29
g30
((lp568
tp569
Rp570
sbatp571
Rp572
sg463
g566
sbsS'Blubb'
p573
g1
(g2
g3
(g173
g573
tp574
tp575
Rp576
(dp577
g9
g423
sg29
g30
((lp578
tp579
Rp580
sbsS'Label'
p581
g1
(g2
g3
(g173
g581
tp582
tp583
Rp584
(dp585
g9
g423
sg29
g30
((lp586
tp587
Rp588
sbsS'Field'
p589
g1
(g2
g3
(g173
g589
tp590
tp591
Rp592
(dp593
g9
g423
sg29
g30
((lp594
tp595
Rp596
sbsS'Exception'
p597
g1
(g2
g3
(g173
g597
tp598
tp599
Rp600
(dp601
g9
g423
sg29
g30
((lp602
tp603
Rp604
sbsS'Namespace'
p605
g1
(g2
g3
(g173
g605
tp606
tp607
Rp608
(dp609
g9
g423
sg29
g30
((lp610
tp611
Rp612
sbsg29
g30
((lp613
g483
ag576
ag521
ag491
ag428
ag600
ag513
ag545
ag561
ag537
ag1
(g2
g3
(g173
g430
tp614
tp615
Rp616
(dp617
g9
g423
sg402
g1
(g2
g3
(g173
g430
g402
tp618
tp619
Rp620
(dp621
g9
g616
sg29
g30
((lp622
tp623
Rp624
sbsg29
g30
((lp625
g1
(g2
g3
(g173
g430
S'Start'
p626
tp627
tp628
Rp629
(dp630
g9
g616
sg29
g30
((lp631
tp632
Rp633
sbag620
atp634
Rp635
sg626
g629
sbag1
(g2
g3
(g173
g57
tp636
tp637
Rp638
(dp639
g9
g423
sS'Member'
p640
g1
(g2
g3
(g173
g57
g640
tp641
tp642
Rp643
(dp644
g9
g638
sg29
g30
((lp645
tp646
Rp647
sbsg29
g30
((lp648
g643
atp649
Rp650
sbag584
ag475
ag608
ag1
(g2
g3
(g173
S'Attribute'
p651
tp652
tp653
Rp654
(dp655
g9
g423
sg425
g1
(g2
g3
(g173
g651
g425
tp656
tp657
Rp658
(dp659
g9
g654
sg29
g30
((lp660
tp661
Rp662
sbsg29
g30
((lp663
g658
atp664
Rp665
sbag553
ag1
(g2
g3
(g173
S'Builtin'
p666
tp667
tp668
Rp669
(dp670
g9
g423
sg526
g1
(g2
g3
(g173
g666
g526
tp671
tp672
Rp673
(dp674
g9
g669
sg29
g30
((lp675
tp676
Rp677
sbsg29
g30
((lp678
g1
(g2
g3
(g173
g666
g518
tp679
tp680
Rp681
(dp682
g9
g669
sg29
g30
((lp683
tp684
Rp685
sbag673
atp686
Rp687
sg518
g681
sbag592
ag529
ag505
atp688
Rp689
sg9
g11
sg430
g616
sg666
g669
sg651
g654
sg57
g638
sbsS'Punctuation'
p690
g1
(g2
g3
(g690
tp691
tp692
Rp693
(dp694
g9
g11
sg29
g30
((lp695
g1
(g2
g3
(g690
S'Indicator'
p696
tp697
tp698
Rp699
(dp700
g9
g693
sg29
g30
((lp701
tp702
Rp703
sbatp704
Rp705
sg696
g699
sbsS'Comment'
p706
g1
(g2
g3
(g706
tp707
tp708
Rp709
(dp710
S'Multi'
p711
g1
(g2
g3
(g706
g711
tp712
tp713
Rp714
(dp715
g9
g709
sg29
g30
((lp716
tp717
Rp718
sbsg9
g11
sS'Special'
p719
g1
(g2
g3
(g706
g719
tp720
tp721
Rp722
(dp723
g9
g709
sg29
g30
((lp724
tp725
Rp726
sbsS'Hashbang'
p727
g1
(g2
g3
(g706
g727
tp728
tp729
Rp730
(dp731
g9
g709
sg29
g30
((lp732
tp733
Rp734
sbsS'Preproc'
p735
g1
(g2
g3
(g706
g735
tp736
tp737
Rp738
(dp739
g9
g709
sg29
g30
((lp740
tp741
Rp742
sbsg214
g1
(g2
g3
(g706
g214
tp743
tp744
Rp745
(dp746
g9
g709
sg29
g30
((lp747
tp748
Rp749
sbsS'Directive'
p750
g1
(g2
g3
(g706
g750
tp751
tp752
Rp753
(dp754
g9
g709
sg29
g30
((lp755
tp756
Rp757
sbsg206
g1
(g2
g3
(g706
g206
tp758
tp759
Rp760
(dp761
g9
g709
sg29
g30
((lp762
tp763
Rp764
sbsS'Singleline'
p765
g1
(g2
g3
(g706
g765
tp766
tp767
Rp768
(dp769
g9
g709
sg29
g30
((lp770
tp771
Rp772
sbsS'Multiline'
p773
g1
(g2
g3
(g706
g773
tp774
tp775
Rp776
(dp777
g9
g709
sg29
g30
((lp778
tp779
Rp780
sbsg29
g30
((lp781
g760
ag753
ag730
ag714
ag768
ag738
ag776
ag745
ag1
(g2
g3
(g706
S'PreprocFile'
p782
tp783
tp784
Rp785
(dp786
g9
g709
sg29
g30
((lp787
tp788
Rp789
sbag1
(g2
g3
(g706
S'SingleLine'
p790
tp791
tp792
Rp793
(dp794
g9
g709
sg29
g30
((lp795
tp796
Rp797
sbag722
atp798
Rp799
sg782
g785
sg790
g793
sbsg14
g39
sg57
g1
(g2
g3
(g57
tp800
tp801
Rp802
(dp803
g9
g11
sg29
g30
((lp804
tp805
Rp806
sbsg370
g1
(g2
g3
(g370
tp807
tp808
Rp809
(dp810
g9
g11
sg29
g30
((lp811
tp812
Rp813
sbsS'Token'
p814
g11
sg197
g1
(g2
g3
(g197
tp815
tp816
Rp817
(dp818
g9
g11
sg29
g30
((lp819
tp820
Rp821
sbsg29
g30
((lp822
g423
ag802
ag7
ag312
ag1
(g2
g3
(S'Text'
p823
tp824
tp825
Rp826
(dp827
S'Beer'
p828
g1
(g2
g3
(g823
g828
tp829
tp830
Rp831
(dp832
g9
g826
sg29
g30
((lp833
tp834
Rp835
sbsS'Whitespace'
p836
g1
(g2
g3
(g823
g836
tp837
tp838
Rp839
(dp840
g9
g826
sg29
g30
((lp841
tp842
Rp843
sbsg9
g11
sS'Root'
p844
g1
(g2
g3
(g823
g844
tp845
tp846
Rp847
(dp848
g9
g826
sg29
g30
((lp849
tp850
Rp851
sbsg101
g1
(g2
g3
(g823
g101
tp852
tp853
Rp854
(dp855
g9
g826
sg29
g30
((lp856
tp857
Rp858
sbsg690
g1
(g2
g3
(g823
g690
tp859
tp860
Rp861
(dp862
g9
g826
sg29
g30
((lp863
tp864
Rp865
sbsg29
g30
((lp866
g847
ag854
ag861
ag839
ag831
ag1
(g2
g3
(g823
S'Rag'
p867
tp868
tp869
Rp870
(dp871
g9
g826
sg29
g30
((lp872
tp873
Rp874
sbatp875
Rp876
sg867
g870
sbag400
ag817
ag693
ag709
ag809
ag39
atp877
Rp878
sg4
g7
sg823
g826
sbsg526
g1
(g2
g3
(g4
g526
tp879
tp880
Rp881
(dp882
g9
g7
sg29
g30
((lp883
tp884
Rp885
sbsS'Control'
p886
g1
(g2
g3
(g4
g886
tp887
tp888
Rp889
(dp890
g9
g7
sg29
g30
((lp891
tp892
Rp893
sbsg550
g1
(g2
g3
(g4
g550
tp894
tp895
Rp896
(dp897
g9
g7
sg29
g30
((lp898
tp899
Rp900
sbsg605
g1
(g2
g3
(g4
g605
tp901
tp902
Rp903
(dp904
g9
g7
sg29
g30
((lp905
tp906
Rp907
sbsS'PreProc'
p908
g1
(g2
g3
(g4
g908
tp909
tp910
Rp911
(dp912
g9
g7
sg29
g30
((lp913
tp914
Rp915
sbsg518
g1
(g2
g3
(g4
g518
tp916
tp917
Rp918
(dp919
g9
g7
sg29
g30
((lp920
tp921
Rp922
sbsS'Reserved'
p923
g1
(g2
g3
(g4
g923
tp924
tp925
Rp926
(dp927
g9
g7
sg29
g30
((lp928
tp929
Rp930
sbsg29
g30
((lp931
g903
ag1
(g2
g3
(g4
g411
tp932
tp933
Rp934
(dp935
g9
g7
sg29
g30
((lp936
tp937
Rp938
sbag889
ag1
(g2
g3
(g4
S'Declaration'
p939
tp940
tp941
Rp942
(dp943
g9
g7
sg29
g30
((lp944
tp945
Rp946
sbag1
(g2
g3
(g4
g4
tp947
tp948
Rp949
(dp950
g9
g7
sg29
g30
((lp951
tp952
Rp953
sbag918
ag896
ag881
ag926
ag911
atp954
Rp955
sg4
g949
sg939
g942
sg411
g934
sbVmodule
p956
tp957
a(g826
V 
p958
tp959
a(g423
Vtoplevel
p960
tp961
a(g693
V(
p962
tp963
a(g423
Vclock
p964
tp965
a(g693
V,
p966
tp967
a(g423
Vreset
p968
tp969
a(g693
V)
p970
tp971
a(g693
V;
p972
tp973
a(g826
V\u000a
p974
tp975
a(g826
g958
tp976
a(g7
Vinput
p977
tp978
a(g826
g958
tp979
a(g423
Vclock
p980
tp981
a(g693
g972
tp982
a(g826
V\u000a
p983
tp984
a(g826
g958
tp985
a(g7
Vinput
p986
tp987
a(g826
g958
tp988
a(g423
Vreset
p989
tp990
a(g693
g972
tp991
a(g826
V\u000a
p992
tp993
a(g826
V \u000a 
p994
tp995
a(g7
Vreg
p996
tp997
a(g826
g958
tp998
a(g423
Vflop1
p999
tp1000
a(g693
g972
tp1001
a(g826
V\u000a
p1002
tp1003
a(g826
g958
tp1004
a(g7
Vreg
p1005
tp1006
a(g826
g958
tp1007
a(g423
Vflop2
p1008
tp1009
a(g693
g972
tp1010
a(g826
V\u000a
p1011
tp1012
a(g826
V \u000a 
p1013
tp1014
a(g7
Valways
p1015
tp1016
a(g826
g958
tp1017
a(g693
V@
p1018
tp1019
a(g826
g958
tp1020
a(g693
g962
tp1021
a(g7
Vposedge
p1022
tp1023
a(g826
g958
tp1024
a(g423
Vreset
p1025
tp1026
a(g826
g958
tp1027
a(g7
Vor
p1028
tp1029
a(g826
g958
tp1030
a(g7
Vposedge
p1031
tp1032
a(g826
g958
tp1033
a(g423
Vclock
p1034
tp1035
a(g693
g970
tp1036
a(g826
V\u000a
p1037
tp1038
a(g826
g958
tp1039
a(g7
Vif
p1040
tp1041
a(g826
g958
tp1042
a(g693
g962
tp1043
a(g423
Vreset
p1044
tp1045
a(g693
g970
tp1046
a(g826
V\u000a
p1047
tp1048
a(g826
V   
p1049
tp1050
a(g7
Vbegin
p1051
tp1052
a(g826
V\u000a
p1053
tp1054
a(g826
V     
p1055
tp1056
a(g423
Vflop1
p1057
tp1058
a(g826
g958
tp1059
a(g400
V<
p1060
tp1061
a(g400
V=
p1062
tp1063
a(g826
g958
tp1064
a(g285
V0
p1065
tp1066
a(g693
g972
tp1067
a(g826
V\u000a
p1068
tp1069
a(g826
V     
p1070
tp1071
a(g423
Vflop2
p1072
tp1073
a(g826
g958
tp1074
a(g400
g1060
tp1075
a(g400
g1062
tp1076
a(g826
g958
tp1077
a(g285
V1
p1078
tp1079
a(g693
g972
tp1080
a(g826
V\u000a
p1081
tp1082
a(g826
V   
p1083
tp1084
a(g7
Vend
p1085
tp1086
a(g826
V\u000a
p1087
tp1088
a(g826
g958
tp1089
a(g7
Velse
p1090
tp1091
a(g826
V\u000a
p1092
tp1093
a(g826
V   
p1094
tp1095
a(g7
Vbegin
p1096
tp1097
a(g826
V\u000a
p1098
tp1099
a(g826
V     
p1100
tp1101
a(g423
Vflop1
p1102
tp1103
a(g826
g958
tp1104
a(g400
g1060
tp1105
a(g400
g1062
tp1106
a(g826
g958
tp1107
a(g423
Vflop2
p1108
tp1109
a(g693
g972
tp1110
a(g826
V\u000a
p1111
tp1112
a(g826
V     
p1113
tp1114
a(g423
Vflop2
p1115
tp1116
a(g826
g958
tp1117
a(g400
g1060
tp1118
a(g400
g1062
tp1119
a(g826
g958
tp1120
a(g423
Vflop1
p1121
tp1122
a(g693
g972
tp1123
a(g826
V\u000a
p1124
tp1125
a(g826
V   
p1126
tp1127
a(g7
Vend
p1128
tp1129
a(g826
V\u000a
p1130
tp1131
a(g7
Vendmodule
p1132
tp1133
a(g826
V\u000a
p1134
tp1135
a.