(lp0
(ccopy_reg
_reconstructor
p1
(cpygments.token
_TokenType
p2
c__builtin__
tuple
p3
(S'Keyword'
p4
tp5
tp6
Rp7
(dp8
S'parent'
p9
g1
(g2
g3
(ttp10
Rp11
(dp12
S'Number'
p13
g1
(g2
g3
(S'Literal'
p14
g13
tp15
tp16
Rp17
(dp18
S'Integer'
p19
g1
(g2
g3
(g14
g13
g19
tp20
tp21
Rp22
(dp23
g9
g17
sS'Long'
p24
g1
(g2
g3
(g14
g13
g19
g24
tp25
tp26
Rp27
(dp28
g9
g22
sS'subtypes'
p29
c__builtin__
set
p30
((lp31
tp32
Rp33
sbsg29
g30
((lp34
g27
atp35
Rp36
sbsg9
g1
(g2
g3
(g14
tp37
tp38
Rp39
(dp40
S'Scalar'
p41
g1
(g2
g3
(g14
g41
tp42
tp43
Rp44
(dp45
g9
g39
sg29
g30
((lp46
g1
(g2
g3
(g14
g41
S'Plain'
p47
tp48
tp49
Rp50
(dp51
g9
g44
sg29
g30
((lp52
tp53
Rp54
sbatp55
Rp56
sg47
g50
sbsg13
g17
sg9
g11
sS'Other'
p57
g1
(g2
g3
(g14
g57
tp58
tp59
Rp60
(dp61
g9
g39
sg29
g30
((lp62
tp63
Rp64
sbsS'Char'
p65
g1
(g2
g3
(g14
g65
tp66
tp67
Rp68
(dp69
g9
g39
sg29
g30
((lp70
tp71
Rp72
sbsS'String'
p73
g1
(g2
g3
(g14
g73
tp74
tp75
Rp76
(dp77
g65
g1
(g2
g3
(g14
g73
g65
tp78
tp79
Rp80
(dp81
g9
g76
sg29
g30
((lp82
tp83
Rp84
sbsS'Backtick'
p85
g1
(g2
g3
(g14
g73
g85
tp86
tp87
Rp88
(dp89
g9
g76
sg29
g30
((lp90
tp91
Rp92
sbsS'Heredoc'
p93
g1
(g2
g3
(g14
g73
g93
tp94
tp95
Rp96
(dp97
g9
g76
sg29
g30
((lp98
tp99
Rp100
sbsS'Symbol'
p101
g1
(g2
g3
(g14
g73
g101
tp102
tp103
Rp104
(dp105
g9
g76
sg29
g30
((lp106
tp107
Rp108
sbsS'Interpol'
p109
g1
(g2
g3
(g14
g73
g109
tp110
tp111
Rp112
(dp113
g9
g76
sg29
g30
((lp114
tp115
Rp116
sbsS'Delimiter'
p117
g1
(g2
g3
(g14
g73
g117
tp118
tp119
Rp120
(dp121
g9
g76
sg29
g30
((lp122
tp123
Rp124
sbsS'Boolean'
p125
g1
(g2
g3
(g14
g73
g125
tp126
tp127
Rp128
(dp129
g9
g76
sg29
g30
((lp130
tp131
Rp132
sbsS'Character'
p133
g1
(g2
g3
(g14
g73
g133
tp134
tp135
Rp136
(dp137
g9
g76
sg29
g30
((lp138
tp139
Rp140
sbsS'Double'
p141
g1
(g2
g3
(g14
g73
g141
tp142
tp143
Rp144
(dp145
g9
g76
sg29
g30
((lp146
tp147
Rp148
sbsS'Delimeter'
p149
g1
(g2
g3
(g14
g73
g149
tp150
tp151
Rp152
(dp153
g9
g76
sg29
g30
((lp154
tp155
Rp156
sbsS'Atom'
p157
g1
(g2
g3
(g14
g73
g157
tp158
tp159
Rp160
(dp161
g9
g76
sg29
g30
((lp162
tp163
Rp164
sbsS'Affix'
p165
g1
(g2
g3
(g14
g73
g165
tp166
tp167
Rp168
(dp169
g9
g76
sg29
g30
((lp170
tp171
Rp172
sbsS'Name'
p173
g1
(g2
g3
(g14
g73
g173
tp174
tp175
Rp176
(dp177
g9
g76
sg29
g30
((lp178
tp179
Rp180
sbsS'Regex'
p181
g1
(g2
g3
(g14
g73
g181
tp182
tp183
Rp184
(dp185
g9
g76
sg29
g30
((lp186
tp187
Rp188
sbsS'Interp'
p189
g1
(g2
g3
(g14
g73
g189
tp190
tp191
Rp192
(dp193
g9
g76
sg29
g30
((lp194
tp195
Rp196
sbsS'Escape'
p197
g1
(g2
g3
(g14
g73
g197
tp198
tp199
Rp200
(dp201
g9
g76
sg29
g30
((lp202
tp203
Rp204
sbsg29
g30
((lp205
g120
ag104
ag184
ag1
(g2
g3
(g14
g73
S'Doc'
p206
tp207
tp208
Rp209
(dp210
g9
g76
sg29
g30
((lp211
tp212
Rp213
sbag136
ag128
ag144
ag112
ag160
ag152
ag176
ag200
ag1
(g2
g3
(g14
g73
S'Single'
p214
tp215
tp216
Rp217
(dp218
g9
g76
sg29
g30
((lp219
tp220
Rp221
sbag1
(g2
g3
(g14
g73
g57
tp222
tp223
Rp224
(dp225
g9
g76
sg29
g30
((lp226
tp227
Rp228
sbag192
ag88
ag168
ag1
(g2
g3
(g14
g73
S'Moment'
p229
tp230
tp231
Rp232
(dp233
g9
g76
sg29
g30
((lp234
tp235
Rp236
sbag80
ag96
atp237
Rp238
sg214
g217
sg229
g232
sg9
g39
sg57
g224
sg206
g209
sbsg29
g30
((lp239
g76
ag68
ag60
ag1
(g2
g3
(g14
S'Date'
p240
tp241
tp242
Rp243
(dp244
g9
g39
sg29
g30
((lp245
tp246
Rp247
sbag44
ag17
atp248
Rp249
sg240
g243
sbsS'Bin'
p250
g1
(g2
g3
(g14
g13
g250
tp251
tp252
Rp253
(dp254
g9
g17
sg29
g30
((lp255
tp256
Rp257
sbsS'Radix'
p258
g1
(g2
g3
(g14
g13
g258
tp259
tp260
Rp261
(dp262
g9
g17
sg29
g30
((lp263
tp264
Rp265
sbsS'Oct'
p266
g1
(g2
g3
(g14
g13
g266
tp267
tp268
Rp269
(dp270
g9
g17
sg29
g30
((lp271
tp272
Rp273
sbsS'Dec'
p274
g1
(g2
g3
(g14
g13
g274
tp275
tp276
Rp277
(dp278
g9
g17
sg29
g30
((lp279
tp280
Rp281
sbsS'Hex'
p282
g1
(g2
g3
(g14
g13
g282
tp283
tp284
Rp285
(dp286
g9
g17
sg29
g30
((lp287
tp288
Rp289
sbsg29
g30
((lp290
g22
ag261
ag277
ag1
(g2
g3
(g14
g13
S'Decimal'
p291
tp292
tp293
Rp294
(dp295
g9
g17
sg29
g30
((lp296
tp297
Rp298
sbag253
ag1
(g2
g3
(g14
g13
S'Float'
p299
tp300
tp301
Rp302
(dp303
g9
g17
sg29
g30
((lp304
tp305
Rp306
sbag269
ag285
atp307
Rp308
sg291
g294
sg299
g302
sbsS'Generic'
p309
g1
(g2
g3
(g309
tp310
tp311
Rp312
(dp313
g9
g11
sS'Deleted'
p314
g1
(g2
g3
(g309
g314
tp315
tp316
Rp317
(dp318
g9
g312
sg29
g30
((lp319
tp320
Rp321
sbsS'Subheading'
p322
g1
(g2
g3
(g309
g322
tp323
tp324
Rp325
(dp326
g9
g312
sg29
g30
((lp327
tp328
Rp329
sbsS'Heading'
p330
g1
(g2
g3
(g309
g330
tp331
tp332
Rp333
(dp334
g9
g312
sg29
g30
((lp335
tp336
Rp337
sbsS'Emph'
p338
g1
(g2
g3
(g309
g338
tp339
tp340
Rp341
(dp342
g9
g312
sg29
g30
((lp343
tp344
Rp345
sbsS'Prompt'
p346
g1
(g2
g3
(g309
g346
tp347
tp348
Rp349
(dp350
g9
g312
sg29
g30
((lp351
tp352
Rp353
sbsS'Inserted'
p354
g1
(g2
g3
(g309
g354
tp355
tp356
Rp357
(dp358
g9
g312
sg29
g30
((lp359
tp360
Rp361
sbsS'Strong'
p362
g1
(g2
g3
(g309
g362
tp363
tp364
Rp365
(dp366
g9
g312
sg29
g30
((lp367
tp368
Rp369
sbsS'Error'
p370
g1
(g2
g3
(g309
g370
tp371
tp372
Rp373
(dp374
g9
g312
sg29
g30
((lp375
tp376
Rp377
sbsS'Traceback'
p378
g1
(g2
g3
(g309
g378
tp379
tp380
Rp381
(dp382
g9
g312
sg29
g30
((lp383
tp384
Rp385
sbsg29
g30
((lp386
g333
ag325
ag1
(g2
g3
(g309
S'Output'
p387
tp388
tp389
Rp390
(dp391
g9
g312
sg29
g30
((lp392
tp393
Rp394
sbag365
ag341
ag373
ag381
ag357
ag349
ag317
atp395
Rp396
sg387
g390
sbsS'Operator'
p397
g1
(g2
g3
(g397
tp398
tp399
Rp400
(dp401
g9
g11
sS'DBS'
p402
g1
(g2
g3
(g397
g402
tp403
tp404
Rp405
(dp406
g9
g400
sg29
g30
((lp407
tp408
Rp409
sbsg29
g30
((lp410
g405
ag1
(g2
g3
(g397
S'Word'
p411
tp412
tp413
Rp414
(dp415
g9
g400
sg29
g30
((lp416
tp417
Rp418
sbatp419
Rp420
sg411
g414
sbsg73
g76
sg173
g1
(g2
g3
(g173
tp421
tp422
Rp423
(dp424
S'Variable'
p425
g1
(g2
g3
(g173
g425
tp426
tp427
Rp428
(dp429
g9
g423
sS'Class'
p430
g1
(g2
g3
(g173
g425
g430
tp431
tp432
Rp433
(dp434
g9
g428
sg29
g30
((lp435
tp436
Rp437
sbsS'Anonymous'
p438
g1
(g2
g3
(g173
g425
g438
tp439
tp440
Rp441
(dp442
g9
g428
sg29
g30
((lp443
tp444
Rp445
sbsS'Instance'
p446
g1
(g2
g3
(g173
g425
g446
tp447
tp448
Rp449
(dp450
g9
g428
sg29
g30
((lp451
tp452
Rp453
sbsS'Global'
p454
g1
(g2
g3
(g173
g425
g454
tp455
tp456
Rp457
(dp458
g9
g428
sg29
g30
((lp459
tp460
Rp461
sbsg29
g30
((lp462
g441
ag449
ag1
(g2
g3
(g173
g425
S'Magic'
p463
tp464
tp465
Rp466
(dp467
g9
g428
sg29
g30
((lp468
tp469
Rp470
sbag457
ag433
atp471
Rp472
sg463
g466
sbsg397
g1
(g2
g3
(g173
g397
tp473
tp474
Rp475
(dp476
g9
g423
sg29
g30
((lp477
tp478
Rp479
sbsS'Decorator'
p480
g1
(g2
g3
(g173
g480
tp481
tp482
Rp483
(dp484
g9
g423
sg29
g30
((lp485
tp486
Rp487
sbsS'Entity'
p488
g1
(g2
g3
(g173
g488
tp489
tp490
Rp491
(dp492
g9
g423
sg402
g1
(g2
g3
(g173
g488
g402
tp493
tp494
Rp495
(dp496
g9
g491
sg29
g30
((lp497
tp498
Rp499
sbsg29
g30
((lp500
g495
atp501
Rp502
sbsg101
g1
(g2
g3
(g173
g101
tp503
tp504
Rp505
(dp506
g9
g423
sg29
g30
((lp507
tp508
Rp509
sbsS'Property'
p510
g1
(g2
g3
(g173
g510
tp511
tp512
Rp513
(dp514
g9
g423
sg29
g30
((lp515
tp516
Rp517
sbsS'Pseudo'
p518
g1
(g2
g3
(g173
g518
tp519
tp520
Rp521
(dp522
g9
g423
sg29
g30
((lp523
tp524
Rp525
sbsS'Type'
p526
g1
(g2
g3
(g173
g526
tp527
tp528
Rp529
(dp530
g9
g423
sg29
g30
((lp531
tp532
Rp533
sbsS'Classes'
p534
g1
(g2
g3
(g173
g534
tp535
tp536
Rp537
(dp538
g9
g423
sg29
g30
((lp539
tp540
Rp541
sbsS'Tag'
p542
g1
(g2
g3
(g173
g542
tp543
tp544
Rp545
(dp546
g9
g423
sg29
g30
((lp547
tp548
Rp549
sbsS'Constant'
p550
g1
(g2
g3
(g173
g550
tp551
tp552
Rp553
(dp554
g9
g423
sg29
g30
((lp555
tp556
Rp557
sbsS'Function'
p558
g1
(g2
g3
(g173
g558
tp559
tp560
Rp561
(dp562
g9
g423
sg29
g30
((lp563
g1
(g2
g3
(g173
g558
g463
tp564
tp565
Rp566
(dp567
g9
g561
sg29
g30
((lp568
tp569
Rp570
sbatp571
Rp572
sg463
g566
sbsS'Blubb'
p573
g1
(g2
g3
(g173
g573
tp574
tp575
Rp576
(dp577
g9
g423
sg29
g30
((lp578
tp579
Rp580
sbsS'Label'
p581
g1
(g2
g3
(g173
g581
tp582
tp583
Rp584
(dp585
g9
g423
sg29
g30
((lp586
tp587
Rp588
sbsS'Field'
p589
g1
(g2
g3
(g173
g589
tp590
tp591
Rp592
(dp593
g9
g423
sg29
g30
((lp594
tp595
Rp596
sbsS'Exception'
p597
g1
(g2
g3
(g173
g597
tp598
tp599
Rp600
(dp601
g9
g423
sg29
g30
((lp602
tp603
Rp604
sbsS'Namespace'
p605
g1
(g2
g3
(g173
g605
tp606
tp607
Rp608
(dp609
g9
g423
sg29
g30
((lp610
tp611
Rp612
sbsg29
g30
((lp613
g483
ag576
ag521
ag491
ag428
ag600
ag513
ag545
ag561
ag537
ag1
(g2
g3
(g173
g430
tp614
tp615
Rp616
(dp617
g9
g423
sg402
g1
(g2
g3
(g173
g430
g402
tp618
tp619
Rp620
(dp621
g9
g616
sg29
g30
((lp622
tp623
Rp624
sbsg29
g30
((lp625
g1
(g2
g3
(g173
g430
S'Start'
p626
tp627
tp628
Rp629
(dp630
g9
g616
sg29
g30
((lp631
tp632
Rp633
sbag620
atp634
Rp635
sg626
g629
sbag1
(g2
g3
(g173
g57
tp636
tp637
Rp638
(dp639
g9
g423
sS'Member'
p640
g1
(g2
g3
(g173
g57
g640
tp641
tp642
Rp643
(dp644
g9
g638
sg29
g30
((lp645
tp646
Rp647
sbsg29
g30
((lp648
g643
atp649
Rp650
sbag584
ag475
ag608
ag1
(g2
g3
(g173
S'Attribute'
p651
tp652
tp653
Rp654
(dp655
g9
g423
sg425
g1
(g2
g3
(g173
g651
g425
tp656
tp657
Rp658
(dp659
g9
g654
sg29
g30
((lp660
tp661
Rp662
sbsg29
g30
((lp663
g658
atp664
Rp665
sbag553
ag1
(g2
g3
(g173
S'Builtin'
p666
tp667
tp668
Rp669
(dp670
g9
g423
sg526
g1
(g2
g3
(g173
g666
g526
tp671
tp672
Rp673
(dp674
g9
g669
sg29
g30
((lp675
tp676
Rp677
sbsg29
g30
((lp678
g1
(g2
g3
(g173
g666
g518
tp679
tp680
Rp681
(dp682
g9
g669
sg29
g30
((lp683
tp684
Rp685
sbag673
atp686
Rp687
sg518
g681
sbag592
ag529
ag505
atp688
Rp689
sg9
g11
sg430
g616
sg666
g669
sg651
g654
sg57
g638
sbsS'Punctuation'
p690
g1
(g2
g3
(g690
tp691
tp692
Rp693
(dp694
g9
g11
sg29
g30
((lp695
g1
(g2
g3
(g690
S'Indicator'
p696
tp697
tp698
Rp699
(dp700
g9
g693
sg29
g30
((lp701
tp702
Rp703
sbatp704
Rp705
sg696
g699
sbsS'Comment'
p706
g1
(g2
g3
(g706
tp707
tp708
Rp709
(dp710
S'Multi'
p711
g1
(g2
g3
(g706
g711
tp712
tp713
Rp714
(dp715
g9
g709
sg29
g30
((lp716
tp717
Rp718
sbsg9
g11
sS'Special'
p719
g1
(g2
g3
(g706
g719
tp720
tp721
Rp722
(dp723
g9
g709
sg29
g30
((lp724
tp725
Rp726
sbsS'Hashbang'
p727
g1
(g2
g3
(g706
g727
tp728
tp729
Rp730
(dp731
g9
g709
sg29
g30
((lp732
tp733
Rp734
sbsS'Preproc'
p735
g1
(g2
g3
(g706
g735
tp736
tp737
Rp738
(dp739
g9
g709
sg29
g30
((lp740
tp741
Rp742
sbsg214
g1
(g2
g3
(g706
g214
tp743
tp744
Rp745
(dp746
g9
g709
sg29
g30
((lp747
tp748
Rp749
sbsS'Directive'
p750
g1
(g2
g3
(g706
g750
tp751
tp752
Rp753
(dp754
g9
g709
sg29
g30
((lp755
tp756
Rp757
sbsg206
g1
(g2
g3
(g706
g206
tp758
tp759
Rp760
(dp761
g9
g709
sg29
g30
((lp762
tp763
Rp764
sbsS'Singleline'
p765
g1
(g2
g3
(g706
g765
tp766
tp767
Rp768
(dp769
g9
g709
sg29
g30
((lp770
tp771
Rp772
sbsS'Multiline'
p773
g1
(g2
g3
(g706
g773
tp774
tp775
Rp776
(dp777
g9
g709
sg29
g30
((lp778
tp779
Rp780
sbsg29
g30
((lp781
g760
ag753
ag730
ag714
ag768
ag738
ag776
ag745
ag1
(g2
g3
(g706
S'PreprocFile'
p782
tp783
tp784
Rp785
(dp786
g9
g709
sg29
g30
((lp787
tp788
Rp789
sbag1
(g2
g3
(g706
S'SingleLine'
p790
tp791
tp792
Rp793
(dp794
g9
g709
sg29
g30
((lp795
tp796
Rp797
sbag722
atp798
Rp799
sg782
g785
sg790
g793
sbsg14
g39
sg57
g1
(g2
g3
(g57
tp800
tp801
Rp802
(dp803
g9
g11
sg29
g30
((lp804
tp805
Rp806
sbsg370
g1
(g2
g3
(g370
tp807
tp808
Rp809
(dp810
g9
g11
sg29
g30
((lp811
tp812
Rp813
sbsS'Token'
p814
g11
sg197
g1
(g2
g3
(g197
tp815
tp816
Rp817
(dp818
g9
g11
sg29
g30
((lp819
tp820
Rp821
sbsg29
g30
((lp822
g423
ag802
ag7
ag312
ag1
(g2
g3
(S'Text'
p823
tp824
tp825
Rp826
(dp827
S'Beer'
p828
g1
(g2
g3
(g823
g828
tp829
tp830
Rp831
(dp832
g9
g826
sg29
g30
((lp833
tp834
Rp835
sbsS'Whitespace'
p836
g1
(g2
g3
(g823
g836
tp837
tp838
Rp839
(dp840
g9
g826
sg29
g30
((lp841
tp842
Rp843
sbsg9
g11
sS'Root'
p844
g1
(g2
g3
(g823
g844
tp845
tp846
Rp847
(dp848
g9
g826
sg29
g30
((lp849
tp850
Rp851
sbsg101
g1
(g2
g3
(g823
g101
tp852
tp853
Rp854
(dp855
g9
g826
sg29
g30
((lp856
tp857
Rp858
sbsg690
g1
(g2
g3
(g823
g690
tp859
tp860
Rp861
(dp862
g9
g826
sg29
g30
((lp863
tp864
Rp865
sbsg29
g30
((lp866
g847
ag854
ag861
ag839
ag831
ag1
(g2
g3
(g823
S'Rag'
p867
tp868
tp869
Rp870
(dp871
g9
g826
sg29
g30
((lp872
tp873
Rp874
sbatp875
Rp876
sg867
g870
sbag400
ag817
ag693
ag709
ag809
ag39
atp877
Rp878
sg4
g7
sg823
g826
sbsg526
g1
(g2
g3
(g4
g526
tp879
tp880
Rp881
(dp882
g9
g7
sg29
g30
((lp883
tp884
Rp885
sbsS'Control'
p886
g1
(g2
g3
(g4
g886
tp887
tp888
Rp889
(dp890
g9
g7
sg29
g30
((lp891
tp892
Rp893
sbsg550
g1
(g2
g3
(g4
g550
tp894
tp895
Rp896
(dp897
g9
g7
sg29
g30
((lp898
tp899
Rp900
sbsg605
g1
(g2
g3
(g4
g605
tp901
tp902
Rp903
(dp904
g9
g7
sg29
g30
((lp905
tp906
Rp907
sbsS'PreProc'
p908
g1
(g2
g3
(g4
g908
tp909
tp910
Rp911
(dp912
g9
g7
sg29
g30
((lp913
tp914
Rp915
sbsg518
g1
(g2
g3
(g4
g518
tp916
tp917
Rp918
(dp919
g9
g7
sg29
g30
((lp920
tp921
Rp922
sbsS'Reserved'
p923
g1
(g2
g3
(g4
g923
tp924
tp925
Rp926
(dp927
g9
g7
sg29
g30
((lp928
tp929
Rp930
sbsg29
g30
((lp931
g903
ag1
(g2
g3
(g4
g411
tp932
tp933
Rp934
(dp935
g9
g7
sg29
g30
((lp936
tp937
Rp938
sbag889
ag1
(g2
g3
(g4
S'Declaration'
p939
tp940
tp941
Rp942
(dp943
g9
g7
sg29
g30
((lp944
tp945
Rp946
sbag1
(g2
g3
(g4
g4
tp947
tp948
Rp949
(dp950
g9
g7
sg29
g30
((lp951
tp952
Rp953
sbag918
ag896
ag881
ag926
ag911
atp954
Rp955
sg4
g949
sg939
g942
sg411
g934
sbVlibrary
p956
tp957
a(g826
V 
p958
tp959
a(g608
Vieee
p960
tp961
a(g693
V;
p962
tp963
a(g826
V\u000a
p964
tp965
a(g7
Vuse
p966
tp967
a(g826
g958
tp968
a(g608
Vieee.std_logic_unsigned.
p969
tp970
a(g7
Vall
p971
tp972
a(g693
g962
tp973
a(g826
V\u000a
p974
tp975
a(g7
Vuse
p976
tp977
a(g826
g958
tp978
a(g608
Vieee.std_logic_1164.
p979
tp980
a(g7
Vall
p981
tp982
a(g693
g962
tp983
a(g826
V   \u000a
p984
tp985
a(g7
Vuse
p986
tp987
a(g826
g958
tp988
a(g608
Vieee.numeric_std.
p989
tp990
a(g7
Vall
p991
tp992
a(g693
g962
tp993
a(g826
V\u000a
p994
tp995
a(g826
V\u000a
p996
tp997
a(g826
V\u000a
p998
tp999
a(g7
Ventity
p1000
tp1001
a(g826
g958
tp1002
a(g616
Vtop_testbench
p1003
tp1004
a(g826
g958
tp1005
a(g7
Vis
p1006
tp1007
a(g826
g958
tp1008
a(g745
V--test
p1009
tp1010
a(g826
V\u000a
p1011
tp1012
a(g826
V	
p1013
tp1014
a(g7
Vgeneric
p1015
tp1016
a(g826
g958
tp1017
a(g693
V(
p1018
tp1019
a(g826
g958
tp1020
a(g745
V-- test
p1021
tp1022
a(g826
V\u000a
p1023
tp1024
a(g826
V	    
p1025
tp1026
a(g423
Vn
p1027
tp1028
a(g826
g958
tp1029
a(g400
V:
p1030
tp1031
a(g826
g958
tp1032
a(g881
Vinteger
p1033
tp1034
a(g826
g958
tp1035
a(g400
g1030
tp1036
a(g400
V=
p1037
tp1038
a(g826
g958
tp1039
a(g22
V8
p1040
tp1041
a(g826
g958
tp1042
a(g745
V-- test
p1043
tp1044
a(g826
V\u000a
p1045
tp1046
a(g826
g1013
tp1047
a(g693
V)
p1048
tp1049
a(g693
g962
tp1050
a(g826
g958
tp1051
a(g745
V-- test
p1052
tp1053
a(g826
V\u000a
p1054
tp1055
a(g7
Vend
p1056
tp1057
a(g826
g958
tp1058
a(g616
Vtop_testbench
p1059
tp1060
a(g693
g962
tp1061
a(g826
g958
tp1062
a(g745
V-- test
p1063
tp1064
a(g826
V\u000a
p1065
tp1066
a(g826
V\u000a
p1067
tp1068
a(g826
V\u000a
p1069
tp1070
a(g7
Varchitecture
p1071
tp1072
a(g826
g958
tp1073
a(g616
Vtop_testbench_arch
p1074
tp1075
a(g826
g958
tp1076
a(g7
Vof
p1077
tp1078
a(g826
g958
tp1079
a(g616
Vtop_testbench
p1080
tp1081
a(g826
g958
tp1082
a(g7
Vis
p1083
tp1084
a(g826
V  \u000a\u000a    
p1085
tp1086
a(g7
Vcomponent
p1087
tp1088
a(g826
g958
tp1089
a(g616
Vtop
p1090
tp1091
a(g826
g958
tp1092
a(g7
Vis
p1093
tp1094
a(g826
V\u000a
p1095
tp1096
a(g826
V        
p1097
tp1098
a(g7
Vgeneric
p1099
tp1100
a(g826
g958
tp1101
a(g693
g1018
tp1102
a(g826
V\u000a
p1103
tp1104
a(g826
V            
p1105
tp1106
a(g423
g1027
tp1107
a(g826
g958
tp1108
a(g400
g1030
tp1109
a(g826
g958
tp1110
a(g881
Vinteger
p1111
tp1112
a(g826
V\u000a
p1113
tp1114
a(g826
V        
p1115
tp1116
a(g693
g1048
tp1117
a(g826
V   
p1118
tp1119
a(g693
g962
tp1120
a(g826
V\u000a
p1121
tp1122
a(g826
V        
p1123
tp1124
a(g7
Vport
p1125
tp1126
a(g826
g958
tp1127
a(g693
g1018
tp1128
a(g826
V\u000a
p1129
tp1130
a(g826
V            
p1131
tp1132
a(g423
Vclk
p1133
tp1134
a(g826
g958
tp1135
a(g400
g1030
tp1136
a(g826
g958
tp1137
a(g7
Vin
p1138
tp1139
a(g826
g958
tp1140
a(g881
Vstd_logic
p1141
tp1142
a(g693
g962
tp1143
a(g826
V\u000a
p1144
tp1145
a(g826
V            
p1146
tp1147
a(g423
Vrst
p1148
tp1149
a(g826
g958
tp1150
a(g400
g1030
tp1151
a(g826
g958
tp1152
a(g7
Vin
p1153
tp1154
a(g826
g958
tp1155
a(g881
Vstd_logic
p1156
tp1157
a(g693
g962
tp1158
a(g826
V\u000a
p1159
tp1160
a(g826
V            
p1161
tp1162
a(g423
Vd1
p1163
tp1164
a(g826
g958
tp1165
a(g400
g1030
tp1166
a(g826
g958
tp1167
a(g7
Vin
p1168
tp1169
a(g826
g958
tp1170
a(g881
Vstd_logic_vector
p1171
tp1172
a(g826
g958
tp1173
a(g693
g1018
tp1174
a(g423
g1027
tp1175
a(g400
V-
p1176
tp1177
a(g22
V1
p1178
tp1179
a(g826
g958
tp1180
a(g7
Vdownto
p1181
tp1182
a(g826
g958
tp1183
a(g22
V0
p1184
tp1185
a(g693
g1048
tp1186
a(g693
g962
tp1187
a(g826
V\u000a
p1188
tp1189
a(g826
V            
p1190
tp1191
a(g423
Vd2
p1192
tp1193
a(g826
g958
tp1194
a(g400
g1030
tp1195
a(g826
g958
tp1196
a(g7
Vin
p1197
tp1198
a(g826
g958
tp1199
a(g881
Vstd_logic_vector
p1200
tp1201
a(g826
g958
tp1202
a(g693
g1018
tp1203
a(g423
g1027
tp1204
a(g400
g1176
tp1205
a(g22
g1178
tp1206
a(g826
g958
tp1207
a(g7
Vdownto
p1208
tp1209
a(g826
g958
tp1210
a(g22
g1184
tp1211
a(g693
g1048
tp1212
a(g693
g962
tp1213
a(g826
V\u000a
p1214
tp1215
a(g826
V            
p1216
tp1217
a(g423
Voperation
p1218
tp1219
a(g826
g958
tp1220
a(g400
g1030
tp1221
a(g826
g958
tp1222
a(g7
Vin
p1223
tp1224
a(g826
g958
tp1225
a(g881
Vstd_logic
p1226
tp1227
a(g693
g962
tp1228
a(g826
V\u000a
p1229
tp1230
a(g826
V            
p1231
tp1232
a(g423
Vresult
p1233
tp1234
a(g826
g958
tp1235
a(g400
g1030
tp1236
a(g826
g958
tp1237
a(g7
Vout
p1238
tp1239
a(g826
g958
tp1240
a(g881
Vstd_logic_vector
p1241
tp1242
a(g826
g958
tp1243
a(g693
g1018
tp1244
a(g22
V2
p1245
tp1246
a(g400
V*
p1247
tp1248
a(g423
g1027
tp1249
a(g400
g1176
tp1250
a(g22
g1178
tp1251
a(g826
g958
tp1252
a(g7
Vdownto
p1253
tp1254
a(g826
g958
tp1255
a(g22
g1184
tp1256
a(g693
g1048
tp1257
a(g826
V\u000a
p1258
tp1259
a(g826
V        
p1260
tp1261
a(g693
g1048
tp1262
a(g693
g962
tp1263
a(g826
V\u000a
p1264
tp1265
a(g826
V    
p1266
tp1267
a(g7
Vend
p1268
tp1269
a(g826
g958
tp1270
a(g7
Vcomponent
p1271
tp1272
a(g693
g962
tp1273
a(g826
V\u000a
p1274
tp1275
a(g826
V\u000a
p1276
tp1277
a(g826
V    
p1278
tp1279
a(g7
Vsignal
p1280
tp1281
a(g826
g958
tp1282
a(g423
Vclk
p1283
tp1284
a(g826
g958
tp1285
a(g400
g1030
tp1286
a(g826
g958
tp1287
a(g881
Vstd_logic
p1288
tp1289
a(g693
g962
tp1290
a(g826
V\u000a
p1291
tp1292
a(g826
V    
p1293
tp1294
a(g7
Vsignal
p1295
tp1296
a(g826
g958
tp1297
a(g423
Vrst
p1298
tp1299
a(g826
g958
tp1300
a(g400
g1030
tp1301
a(g826
g958
tp1302
a(g881
Vstd_logic
p1303
tp1304
a(g693
g962
tp1305
a(g826
V\u000a
p1306
tp1307
a(g826
g1013
tp1308
a(g7
Vsignal
p1309
tp1310
a(g826
g958
tp1311
a(g423
Voperation
p1312
tp1313
a(g826
g958
tp1314
a(g400
g1030
tp1315
a(g826
g958
tp1316
a(g881
Vstd_logic
p1317
tp1318
a(g693
g962
tp1319
a(g826
V\u000a
p1320
tp1321
a(g826
V    
p1322
tp1323
a(g7
Vsignal
p1324
tp1325
a(g826
g958
tp1326
a(g423
Vd1
p1327
tp1328
a(g826
g958
tp1329
a(g400
g1030
tp1330
a(g826
g958
tp1331
a(g881
Vstd_logic_vector
p1332
tp1333
a(g826
g958
tp1334
a(g693
g1018
tp1335
a(g423
g1027
tp1336
a(g400
g1176
tp1337
a(g22
g1178
tp1338
a(g826
g958
tp1339
a(g7
Vdownto
p1340
tp1341
a(g826
g958
tp1342
a(g22
g1184
tp1343
a(g693
g1048
tp1344
a(g693
g962
tp1345
a(g826
V\u000a
p1346
tp1347
a(g826
V    
p1348
tp1349
a(g7
Vsignal
p1350
tp1351
a(g826
g958
tp1352
a(g423
Vd2
p1353
tp1354
a(g826
g958
tp1355
a(g400
g1030
tp1356
a(g826
g958
tp1357
a(g881
Vstd_logic_vector
p1358
tp1359
a(g826
g958
tp1360
a(g693
g1018
tp1361
a(g423
g1027
tp1362
a(g400
g1176
tp1363
a(g22
g1178
tp1364
a(g826
g958
tp1365
a(g7
Vdownto
p1366
tp1367
a(g826
g958
tp1368
a(g22
g1184
tp1369
a(g693
g1048
tp1370
a(g693
g962
tp1371
a(g826
V\u000a
p1372
tp1373
a(g826
V    
p1374
tp1375
a(g7
Vsignal
p1376
tp1377
a(g826
g958
tp1378
a(g423
Vresult
p1379
tp1380
a(g826
g958
tp1381
a(g400
g1030
tp1382
a(g826
g958
tp1383
a(g881
Vstd_logic_vector
p1384
tp1385
a(g826
g958
tp1386
a(g693
g1018
tp1387
a(g22
g1245
tp1388
a(g400
g1247
tp1389
a(g423
g1027
tp1390
a(g400
g1176
tp1391
a(g22
g1178
tp1392
a(g826
g958
tp1393
a(g7
Vdownto
p1394
tp1395
a(g826
g958
tp1396
a(g22
g1184
tp1397
a(g693
g1048
tp1398
a(g693
g962
tp1399
a(g826
V\u000a
p1400
tp1401
a(g826
V    \u000a    
p1402
tp1403
a(g7
Vtype
p1404
tp1405
a(g826
g958
tp1406
a(g423
Vtest_type
p1407
tp1408
a(g826
g958
tp1409
a(g7
Vis
p1410
tp1411
a(g826
g958
tp1412
a(g693
g1018
tp1413
a(g826
g958
tp1414
a(g423
Va1
p1415
tp1416
a(g693
V,
p1417
tp1418
a(g826
g958
tp1419
a(g423
Va2
p1420
tp1421
a(g693
g1417
tp1422
a(g826
g958
tp1423
a(g423
Va3
p1424
tp1425
a(g693
g1417
tp1426
a(g826
g958
tp1427
a(g423
Va4
p1428
tp1429
a(g693
g1417
tp1430
a(g826
g958
tp1431
a(g423
Va5
p1432
tp1433
a(g693
g1417
tp1434
a(g826
g958
tp1435
a(g423
Va6
p1436
tp1437
a(g693
g1417
tp1438
a(g826
g958
tp1439
a(g423
Va7
p1440
tp1441
a(g693
g1417
tp1442
a(g826
g958
tp1443
a(g423
Va8
p1444
tp1445
a(g693
g1417
tp1446
a(g826
g958
tp1447
a(g423
Va9
p1448
tp1449
a(g693
g1417
tp1450
a(g826
g958
tp1451
a(g423
Va10
p1452
tp1453
a(g693
g1048
tp1454
a(g693
g962
tp1455
a(g826
V\u000a
p1456
tp1457
a(g826
V    
p1458
tp1459
a(g7
Vattribute
p1460
tp1461
a(g826
g958
tp1462
a(g423
Venum_encoding
p1463
tp1464
a(g826
g958
tp1465
a(g7
Vof
p1466
tp1467
a(g826
g958
tp1468
a(g423
Vmy_state
p1469
tp1470
a(g826
g958
tp1471
a(g400
g1030
tp1472
a(g826
g958
tp1473
a(g7
Vtype
p1474
tp1475
a(g826
g958
tp1476
a(g7
Vis
p1477
tp1478
a(g826
g958
tp1479
a(g76
V"001 010 011 100 111"
p1480
tp1481
a(g693
g962
tp1482
a(g826
V\u000a
p1483
tp1484
a(g7
Vbegin
p1485
tp1486
a(g826
V\u000a
p1487
tp1488
a(g826
V\u000a
p1489
tp1490
a(g826
V    
p1491
tp1492
a(g423
VTESTUNIT
p1493
tp1494
a(g826
g958
tp1495
a(g400
g1030
tp1496
a(g826
g958
tp1497
a(g423
Vtop
p1498
tp1499
a(g826
g958
tp1500
a(g7
Vgeneric
p1501
tp1502
a(g826
g958
tp1503
a(g7
Vmap
p1504
tp1505
a(g826
g958
tp1506
a(g693
g1018
tp1507
a(g423
g1027
tp1508
a(g826
g958
tp1509
a(g400
g1037
tp1510
a(g400
V>
p1511
tp1512
a(g826
g958
tp1513
a(g423
g1027
tp1514
a(g693
g1048
tp1515
a(g826
V\u000a
p1516
tp1517
a(g826
V                   
p1518
tp1519
a(g7
Vport
p1520
tp1521
a(g826
g958
tp1522
a(g7
Vmap
p1523
tp1524
a(g826
g958
tp1525
a(g693
g1018
tp1526
a(g423
Vclk
p1527
tp1528
a(g826
g958
tp1529
a(g400
g1037
tp1530
a(g400
g1511
tp1531
a(g826
g958
tp1532
a(g423
Vclk
p1533
tp1534
a(g693
g1417
tp1535
a(g826
V\u000a
p1536
tp1537
a(g826
V                             
p1538
tp1539
a(g423
Vrst
p1540
tp1541
a(g826
g958
tp1542
a(g400
g1037
tp1543
a(g400
g1511
tp1544
a(g826
g958
tp1545
a(g423
Vrst
p1546
tp1547
a(g693
g1417
tp1548
a(g826
V\u000a
p1549
tp1550
a(g826
V                             
p1551
tp1552
a(g423
Vd1
p1553
tp1554
a(g826
V  
p1555
tp1556
a(g400
g1037
tp1557
a(g400
g1511
tp1558
a(g826
g958
tp1559
a(g423
Vd1
p1560
tp1561
a(g693
g1417
tp1562
a(g826
V\u000a
p1563
tp1564
a(g826
V                             
p1565
tp1566
a(g423
Vd2
p1567
tp1568
a(g826
V  
p1569
tp1570
a(g400
g1037
tp1571
a(g400
g1511
tp1572
a(g826
g958
tp1573
a(g423
Vd2
p1574
tp1575
a(g693
g1417
tp1576
a(g826
V\u000a
p1577
tp1578
a(g826
V                             
p1579
tp1580
a(g423
Voperation
p1581
tp1582
a(g826
g958
tp1583
a(g400
g1037
tp1584
a(g400
g1511
tp1585
a(g826
g958
tp1586
a(g423
Voperation
p1587
tp1588
a(g693
g1417
tp1589
a(g826
V\u000a
p1590
tp1591
a(g826
V                             
p1592
tp1593
a(g423
Vresult
p1594
tp1595
a(g826
g958
tp1596
a(g400
g1037
tp1597
a(g400
g1511
tp1598
a(g826
g958
tp1599
a(g423
Vresult
p1600
tp1601
a(g693
g1048
tp1602
a(g693
g962
tp1603
a(g826
V\u000a
p1604
tp1605
a(g826
V\u000a
p1606
tp1607
a(g826
V    
p1608
tp1609
a(g423
Vclock_process
p1610
tp1611
a(g826
g958
tp1612
a(g400
g1030
tp1613
a(g826
g958
tp1614
a(g7
Vprocess
p1615
tp1616
a(g826
V\u000a
p1617
tp1618
a(g826
V    
p1619
tp1620
a(g7
Vbegin
p1621
tp1622
a(g826
V\u000a
p1623
tp1624
a(g826
V        
p1625
tp1626
a(g423
Vclk
p1627
tp1628
a(g826
g958
tp1629
a(g400
V<
p1630
tp1631
a(g400
g1037
tp1632
a(g826
g958
tp1633
a(g80
V'0'
p1634
tp1635
a(g693
g962
tp1636
a(g826
V\u000a
p1637
tp1638
a(g826
V        
p1639
tp1640
a(g7
Vwait
p1641
tp1642
a(g826
g958
tp1643
a(g7
Vfor
p1644
tp1645
a(g826
g958
tp1646
a(g22
V5
p1647
tp1648
a(g826
g958
tp1649
a(g423
Vns
p1650
tp1651
a(g693
g962
tp1652
a(g826
V\u000a
p1653
tp1654
a(g826
V        
p1655
tp1656
a(g423
Vclk
p1657
tp1658
a(g826
g958
tp1659
a(g400
g1630
tp1660
a(g400
g1037
tp1661
a(g826
g958
tp1662
a(g80
V'1'
p1663
tp1664
a(g693
g962
tp1665
a(g826
V\u000a
p1666
tp1667
a(g826
V        
p1668
tp1669
a(g7
Vwait
p1670
tp1671
a(g826
g958
tp1672
a(g7
Vfor
p1673
tp1674
a(g826
g958
tp1675
a(g22
g1647
tp1676
a(g826
g958
tp1677
a(g423
Vns
p1678
tp1679
a(g693
g962
tp1680
a(g826
V\u000a
p1681
tp1682
a(g826
V    
p1683
tp1684
a(g7
Vend
p1685
tp1686
a(g826
g958
tp1687
a(g7
Vprocess
p1688
tp1689
a(g693
g962
tp1690
a(g826
V\u000a
p1691
tp1692
a(g826
V\u000a
p1693
tp1694
a(g826
V    
p1695
tp1696
a(g423
Vdata_process
p1697
tp1698
a(g826
g958
tp1699
a(g400
g1030
tp1700
a(g826
g958
tp1701
a(g7
Vprocess
p1702
tp1703
a(g826
V\u000a
p1704
tp1705
a(g826
V    
p1706
tp1707
a(g7
Vbegin
p1708
tp1709
a(g826
V       \u000a		\u000a		
p1710
tp1711
a(g745
V-- test case #1	
p1712
tp1713
a(g826
V\u000a
p1714
tp1715
a(g826
V	   	
p1716
tp1717
a(g423
Voperation
p1718
tp1719
a(g826
g958
tp1720
a(g400
g1630
tp1721
a(g400
g1037
tp1722
a(g826
g958
tp1723
a(g80
V'0'
p1724
tp1725
a(g693
g962
tp1726
a(g826
V\u000a
p1727
tp1728
a(g826
V		\u000a        
p1729
tp1730
a(g423
Vrst
p1731
tp1732
a(g826
g958
tp1733
a(g400
g1630
tp1734
a(g400
g1037
tp1735
a(g826
g958
tp1736
a(g80
V'1'
p1737
tp1738
a(g693
g962
tp1739
a(g826
V\u000a
p1740
tp1741
a(g826
V        
p1742
tp1743
a(g7
Vwait
p1744
tp1745
a(g826
g958
tp1746
a(g7
Vfor
p1747
tp1748
a(g826
g958
tp1749
a(g22
g1647
tp1750
a(g826
g958
tp1751
a(g423
Vns
p1752
tp1753
a(g693
g962
tp1754
a(g826
V\u000a
p1755
tp1756
a(g826
V        
p1757
tp1758
a(g423
Vrst
p1759
tp1760
a(g826
g958
tp1761
a(g400
g1630
tp1762
a(g400
g1037
tp1763
a(g826
g958
tp1764
a(g80
V'0'
p1765
tp1766
a(g693
g962
tp1767
a(g826
V\u000a
p1768
tp1769
a(g826
V        
p1770
tp1771
a(g7
Vwait
p1772
tp1773
a(g826
g958
tp1774
a(g7
Vfor
p1775
tp1776
a(g826
g958
tp1777
a(g22
g1647
tp1778
a(g826
g958
tp1779
a(g423
Vns
p1780
tp1781
a(g693
g962
tp1782
a(g826
V\u000a
p1783
tp1784
a(g826
V		\u000a		
p1785
tp1786
a(g423
Vd1
p1787
tp1788
a(g826
g958
tp1789
a(g400
g1630
tp1790
a(g400
g1037
tp1791
a(g826
g958
tp1792
a(g881
Vstd_logic_vector
p1793
tp1794
a(g693
g1018
tp1795
a(g423
Vto_unsigned
p1796
tp1797
a(g693
g1018
tp1798
a(g22
V60
p1799
tp1800
a(g693
g1417
tp1801
a(g826
g958
tp1802
a(g423
Vd1
p1803
tp1804
a(g654
V'length
p1805
tp1806
a(g693
g1048
tp1807
a(g693
g1048
tp1808
a(g693
g962
tp1809
a(g826
V\u000a
p1810
tp1811
a(g826
V		
p1812
tp1813
a(g423
Vd2
p1814
tp1815
a(g826
g958
tp1816
a(g400
g1630
tp1817
a(g400
g1037
tp1818
a(g826
g958
tp1819
a(g881
Vstd_logic_vector
p1820
tp1821
a(g693
g1018
tp1822
a(g423
Vto_unsigned
p1823
tp1824
a(g693
g1018
tp1825
a(g22
V12
p1826
tp1827
a(g693
g1417
tp1828
a(g826
g958
tp1829
a(g423
Vd2
p1830
tp1831
a(g654
V'length
p1832
tp1833
a(g693
g1048
tp1834
a(g693
g1048
tp1835
a(g693
g962
tp1836
a(g826
V\u000a
p1837
tp1838
a(g826
V		
p1839
tp1840
a(g7
Vwait
p1841
tp1842
a(g826
g958
tp1843
a(g7
Vfor
p1844
tp1845
a(g826
g958
tp1846
a(g22
V360
p1847
tp1848
a(g826
g958
tp1849
a(g423
Vns
p1850
tp1851
a(g693
g962
tp1852
a(g826
V\u000a
p1853
tp1854
a(g826
V		\u000a		
p1855
tp1856
a(g7
Vassert
p1857
tp1858
a(g826
g958
tp1859
a(g693
g1018
tp1860
a(g423
Vresult
p1861
tp1862
a(g826
g958
tp1863
a(g400
g1037
tp1864
a(g826
g958
tp1865
a(g881
Vstd_logic_vector
p1866
tp1867
a(g693
g1018
tp1868
a(g423
Vto_unsigned
p1869
tp1870
a(g693
g1018
tp1871
a(g22
V720
p1872
tp1873
a(g693
g1417
tp1874
a(g826
g958
tp1875
a(g423
Vresult
p1876
tp1877
a(g654
V'length
p1878
tp1879
a(g693
g1048
tp1880
a(g693
g1048
tp1881
a(g693
g1048
tp1882
a(g826
V\u000a
p1883
tp1884
a(g826
V			
p1885
tp1886
a(g423
Vreport
p1887
tp1888
a(g826
g958
tp1889
a(g76
V"Test case #1 failed"
p1890
tp1891
a(g826
g958
tp1892
a(g7
Vseverity
p1893
tp1894
a(g826
g958
tp1895
a(g423
Verror
p1896
tp1897
a(g693
g962
tp1898
a(g826
V \u000a            \u000a		
p1899
tp1900
a(g745
V-- test case #2	
p1901
tp1902
a(g826
V\u000a
p1903
tp1904
a(g826
V	   	
p1905
tp1906
a(g423
Voperation
p1907
tp1908
a(g826
g958
tp1909
a(g400
g1630
tp1910
a(g400
g1037
tp1911
a(g826
g958
tp1912
a(g80
V'0'
p1913
tp1914
a(g693
g962
tp1915
a(g826
V\u000a
p1916
tp1917
a(g826
V		\u000a        
p1918
tp1919
a(g423
Vrst
p1920
tp1921
a(g826
g958
tp1922
a(g400
g1630
tp1923
a(g400
g1037
tp1924
a(g826
g958
tp1925
a(g80
V'1'
p1926
tp1927
a(g693
g962
tp1928
a(g826
V\u000a
p1929
tp1930
a(g826
V        
p1931
tp1932
a(g7
Vwait
p1933
tp1934
a(g826
g958
tp1935
a(g7
Vfor
p1936
tp1937
a(g826
g958
tp1938
a(g22
g1647
tp1939
a(g826
g958
tp1940
a(g423
Vns
p1941
tp1942
a(g693
g962
tp1943
a(g826
V\u000a
p1944
tp1945
a(g826
V        
p1946
tp1947
a(g423
Vrst
p1948
tp1949
a(g826
g958
tp1950
a(g400
g1630
tp1951
a(g400
g1037
tp1952
a(g826
g958
tp1953
a(g80
V'0'
p1954
tp1955
a(g693
g962
tp1956
a(g826
V\u000a
p1957
tp1958
a(g826
V        
p1959
tp1960
a(g7
Vwait
p1961
tp1962
a(g826
g958
tp1963
a(g7
Vfor
p1964
tp1965
a(g826
g958
tp1966
a(g22
g1647
tp1967
a(g826
g958
tp1968
a(g423
Vns
p1969
tp1970
a(g693
g962
tp1971
a(g826
V\u000a
p1972
tp1973
a(g826
V		\u000a		
p1974
tp1975
a(g423
Vd1
p1976
tp1977
a(g826
g958
tp1978
a(g400
g1630
tp1979
a(g400
g1037
tp1980
a(g826
g958
tp1981
a(g881
Vstd_logic_vector
p1982
tp1983
a(g693
g1018
tp1984
a(g423
Vto_unsigned
p1985
tp1986
a(g693
g1018
tp1987
a(g22
V55
p1988
tp1989
a(g693
g1417
tp1990
a(g826
g958
tp1991
a(g423
Vd1
p1992
tp1993
a(g654
V'length
p1994
tp1995
a(g693
g1048
tp1996
a(g693
g1048
tp1997
a(g693
g962
tp1998
a(g826
V\u000a
p1999
tp2000
a(g826
V		
p2001
tp2002
a(g423
Vd2
p2003
tp2004
a(g826
g958
tp2005
a(g400
g1630
tp2006
a(g400
g1037
tp2007
a(g826
g958
tp2008
a(g881
Vstd_logic_vector
p2009
tp2010
a(g693
g1018
tp2011
a(g423
Vto_unsigned
p2012
tp2013
a(g693
g1018
tp2014
a(g22
g1178
tp2015
a(g693
g1417
tp2016
a(g826
g958
tp2017
a(g423
Vd2
p2018
tp2019
a(g654
V'length
p2020
tp2021
a(g693
g1048
tp2022
a(g693
g1048
tp2023
a(g693
g962
tp2024
a(g826
V\u000a
p2025
tp2026
a(g826
V		
p2027
tp2028
a(g7
Vwait
p2029
tp2030
a(g826
g958
tp2031
a(g7
Vfor
p2032
tp2033
a(g826
g958
tp2034
a(g22
V360
p2035
tp2036
a(g826
g958
tp2037
a(g423
Vns
p2038
tp2039
a(g693
g962
tp2040
a(g826
V\u000a
p2041
tp2042
a(g826
V		\u000a		
p2043
tp2044
a(g7
Vassert
p2045
tp2046
a(g826
g958
tp2047
a(g693
g1018
tp2048
a(g423
Vresult
p2049
tp2050
a(g826
g958
tp2051
a(g400
g1037
tp2052
a(g826
g958
tp2053
a(g881
Vstd_logic_vector
p2054
tp2055
a(g693
g1018
tp2056
a(g423
Vto_unsigned
p2057
tp2058
a(g693
g1018
tp2059
a(g22
V55
p2060
tp2061
a(g693
g1417
tp2062
a(g826
g958
tp2063
a(g423
Vresult
p2064
tp2065
a(g654
V'length
p2066
tp2067
a(g693
g1048
tp2068
a(g693
g1048
tp2069
a(g693
g1048
tp2070
a(g826
V\u000a
p2071
tp2072
a(g826
V			
p2073
tp2074
a(g423
Vreport
p2075
tp2076
a(g826
g958
tp2077
a(g76
V"Test case #2 failed"
p2078
tp2079
a(g826
g958
tp2080
a(g7
Vseverity
p2081
tp2082
a(g826
g958
tp2083
a(g423
Verror
p2084
tp2085
a(g693
g962
tp2086
a(g826
V\u000a
p2087
tp2088
a(g826
V            \u000a        
p2089
tp2090
a(g745
V-- etc 
p2091
tp2092
a(g826
V\u000a
p2093
tp2094
a(g826
V            \u000a    
p2095
tp2096
a(g7
Vend
p2097
tp2098
a(g826
g958
tp2099
a(g7
Vprocess
p2100
tp2101
a(g693
g962
tp2102
a(g826
V\u000a
p2103
tp2104
a(g826
V\u000a
p2105
tp2106
a(g7
Vend
p2107
tp2108
a(g826
g958
tp2109
a(g616
Vtop_testbench_arch
p2110
tp2111
a(g693
g962
tp2112
a(g826
V\u000a
p2113
tp2114
a(g826
V\u000a
p2115
tp2116
a(g826
V\u000a
p2117
tp2118
a(g7
Vconfiguration
p2119
tp2120
a(g826
g958
tp2121
a(g616
Vtestbench_for_top
p2122
tp2123
a(g826
g958
tp2124
a(g7
Vof
p2125
tp2126
a(g826
g958
tp2127
a(g616
Vtop_testbench
p2128
tp2129
a(g826
g958
tp2130
a(g7
Vis
p2131
tp2132
a(g826
V\u000a
p2133
tp2134
a(g826
g1013
tp2135
a(g7
Vfor
p2136
tp2137
a(g826
g958
tp2138
a(g423
Vtop_testbench_arch
p2139
tp2140
a(g826
V\u000a
p2141
tp2142
a(g826
V		
p2143
tp2144
a(g7
Vfor
p2145
tp2146
a(g826
g958
tp2147
a(g423
VTESTUNIT
p2148
tp2149
a(g826
g958
tp2150
a(g400
g1030
tp2151
a(g826
g958
tp2152
a(g423
Vtop
p2153
tp2154
a(g826
V\u000a
p2155
tp2156
a(g826
V			
p2157
tp2158
a(g7
Vuse
p2159
tp2160
a(g826
g958
tp2161
a(g7
Ventity
p2162
tp2163
a(g826
g958
tp2164
a(g608
Vwork
p2165
tp2166
a(g693
V.
p2167
tp2168
a(g423
Vtop
p2169
tp2170
a(g693
g1018
tp2171
a(g423
Vtop_arch
p2172
tp2173
a(g693
g1048
tp2174
a(g693
g962
tp2175
a(g826
V\u000a
p2176
tp2177
a(g826
V		
p2178
tp2179
a(g7
Vend
p2180
tp2181
a(g826
g958
tp2182
a(g7
Vfor
p2183
tp2184
a(g693
g962
tp2185
a(g826
V\u000a
p2186
tp2187
a(g826
g1013
tp2188
a(g7
Vend
p2189
tp2190
a(g826
g958
tp2191
a(g7
Vfor
p2192
tp2193
a(g693
g962
tp2194
a(g826
V\u000a
p2195
tp2196
a(g7
Vend
p2197
tp2198
a(g826
g958
tp2199
a(g616
Vtestbench_for_top
p2200
tp2201
a(g693
g962
tp2202
a(g826
V\u000a
p2203
tp2204
a(g826
V\u000a
p2205
tp2206
a(g826
V\u000a
p2207
tp2208
a(g7
Vfunction
p2209
tp2210
a(g826
g958
tp2211
a(g423
Vcompare
p2212
tp2213
a(g693
g1018
tp2214
a(g423
VA
p2215
tp2216
a(g400
g1030
tp2217
a(g826
g958
tp2218
a(g881
Vstd_logic
p2219
tp2220
a(g693
g1417
tp2221
a(g826
g958
tp2222
a(g423
VB
p2223
tp2224
a(g400
g1030
tp2225
a(g826
g958
tp2226
a(g881
Vstd_Logic
p2227
tp2228
a(g693
g1048
tp2229
a(g826
g958
tp2230
a(g7
Vreturn
p2231
tp2232
a(g826
g958
tp2233
a(g881
Vstd_logic
p2234
tp2235
a(g826
g958
tp2236
a(g7
Vis
p2237
tp2238
a(g826
V\u000a
p2239
tp2240
a(g826
V    
p2241
tp2242
a(g7
Vconstant
p2243
tp2244
a(g826
g958
tp2245
a(g423
Vpi
p2246
tp2247
a(g826
g958
tp2248
a(g400
g1030
tp2249
a(g826
g958
tp2250
a(g423
Vreal
p2251
tp2252
a(g826
g958
tp2253
a(g400
g1030
tp2254
a(g400
g1037
tp2255
a(g826
g958
tp2256
a(g22
V3
p2257
tp2258
a(g693
g2167
tp2259
a(g22
V14159
p2260
tp2261
a(g693
g962
tp2262
a(g826
V\u000a
p2263
tp2264
a(g826
V    
p2265
tp2266
a(g7
Vconstant
p2267
tp2268
a(g826
g958
tp2269
a(g423
Vhalf_pi
p2270
tp2271
a(g826
g958
tp2272
a(g400
g1030
tp2273
a(g826
g958
tp2274
a(g423
Vreal
p2275
tp2276
a(g826
g958
tp2277
a(g400
g1030
tp2278
a(g400
g1037
tp2279
a(g826
g958
tp2280
a(g423
Vpi
p2281
tp2282
a(g826
g958
tp2283
a(g400
V/
p2284
tp2285
a(g826
g958
tp2286
a(g22
g1245
tp2287
a(g693
g2167
tp2288
a(g22
g1184
tp2289
a(g693
g962
tp2290
a(g826
V\u000a
p2291
tp2292
a(g826
V    
p2293
tp2294
a(g7
Vconstant
p2295
tp2296
a(g826
g958
tp2297
a(g423
Vcycle_time
p2298
tp2299
a(g826
g958
tp2300
a(g400
g1030
tp2301
a(g826
g958
tp2302
a(g881
Vtime
p2303
tp2304
a(g826
g958
tp2305
a(g400
g1030
tp2306
a(g400
g1037
tp2307
a(g826
g958
tp2308
a(g22
g1245
tp2309
a(g826
g958
tp2310
a(g423
Vns
p2311
tp2312
a(g693
g962
tp2313
a(g826
V\u000a
p2314
tp2315
a(g826
V    
p2316
tp2317
a(g7
Vconstant
p2318
tp2319
a(g826
g958
tp2320
a(g423
VN
p2321
tp2322
a(g693
g1417
tp2323
a(g826
g958
tp2324
a(g423
VN5
p2325
tp2326
a(g826
g958
tp2327
a(g400
g1030
tp2328
a(g826
g958
tp2329
a(g881
Vinteger
p2330
tp2331
a(g826
g958
tp2332
a(g400
g1030
tp2333
a(g400
g1037
tp2334
a(g826
g958
tp2335
a(g22
g1647
tp2336
a(g693
g962
tp2337
a(g826
V\u000a
p2338
tp2339
a(g7
Vbegin
p2340
tp2341
a(g826
V\u000a
p2342
tp2343
a(g826
V    
p2344
tp2345
a(g7
Vif
p2346
tp2347
a(g826
g958
tp2348
a(g693
g1018
tp2349
a(g423
g2215
tp2350
a(g826
g958
tp2351
a(g400
g1037
tp2352
a(g826
g958
tp2353
a(g80
V'0'
p2354
tp2355
a(g826
g958
tp2356
a(g7
Vand
p2357
tp2358
a(g826
g958
tp2359
a(g423
g2223
tp2360
a(g826
g958
tp2361
a(g400
g1037
tp2362
a(g826
g958
tp2363
a(g80
V'1'
p2364
tp2365
a(g693
g1048
tp2366
a(g826
g958
tp2367
a(g7
Vthen
p2368
tp2369
a(g826
V\u000a
p2370
tp2371
a(g826
V        
p2372
tp2373
a(g7
Vreturn
p2374
tp2375
a(g826
g958
tp2376
a(g423
g2223
tp2377
a(g693
g962
tp2378
a(g826
V\u000a
p2379
tp2380
a(g826
V    
p2381
tp2382
a(g7
Velse
p2383
tp2384
a(g826
V\u000a
p2385
tp2386
a(g826
V        
p2387
tp2388
a(g7
Vreturn
p2389
tp2390
a(g826
g958
tp2391
a(g423
g2215
tp2392
a(g693
g962
tp2393
a(g826
V\u000a
p2394
tp2395
a(g826
V    
p2396
tp2397
a(g7
Vend
p2398
tp2399
a(g826
g958
tp2400
a(g7
Vif
p2401
tp2402
a(g826
g958
tp2403
a(g693
g962
tp2404
a(g826
V\u000a
p2405
tp2406
a(g7
Vend
p2407
tp2408
a(g826
g958
tp2409
a(g616
Vcompare
p2410
tp2411
a(g693
g962
tp2412
a(g826
V\u000a
p2413
tp2414
a(g826
V\u000a
p2415
tp2416
a(g826
V\u000a
p2417
tp2418
a(g7
Vprocedure
p2419
tp2420
a(g826
g958
tp2421
a(g423
Vprint
p2422
tp2423
a(g693
g1018
tp2424
a(g423
VP
p2425
tp2426
a(g826
g958
tp2427
a(g400
g1030
tp2428
a(g826
g958
tp2429
a(g881
Vstd_logic_vector
p2430
tp2431
a(g693
g1018
tp2432
a(g22
V7
p2433
tp2434
a(g826
g958
tp2435
a(g7
Vdownto
p2436
tp2437
a(g826
g958
tp2438
a(g22
g1184
tp2439
a(g693
g1048
tp2440
a(g693
g962
tp2441
a(g826
V\u000a
p2442
tp2443
a(g826
V                
p2444
tp2445
a(g423
VU
p2446
tp2447
a(g826
g958
tp2448
a(g400
g1030
tp2449
a(g826
g958
tp2450
a(g881
Vstd_logic_vector
p2451
tp2452
a(g693
g1018
tp2453
a(g22
g2257
tp2454
a(g826
g958
tp2455
a(g7
Vdownto
p2456
tp2457
a(g826
g958
tp2458
a(g22
g1184
tp2459
a(g693
g1048
tp2460
a(g693
g1048
tp2461
a(g826
g958
tp2462
a(g7
Vis
p2463
tp2464
a(g826
V\u000a
p2465
tp2466
a(g826
V    
p2467
tp2468
a(g7
Vvariable
p2469
tp2470
a(g826
g958
tp2471
a(g423
Vmy_line
p2472
tp2473
a(g826
g958
tp2474
a(g400
g1030
tp2475
a(g826
g958
tp2476
a(g423
Vline
p2477
tp2478
a(g693
g962
tp2479
a(g826
V\u000a
p2480
tp2481
a(g826
V    
p2482
tp2483
a(g7
Valias
p2484
tp2485
a(g826
g958
tp2486
a(g423
Vswrite
p2487
tp2488
a(g826
g958
tp2489
a(g7
Vis
p2490
tp2491
a(g826
g958
tp2492
a(g423
Vwrite
p2493
tp2494
a(g826
g958
tp2495
a(g693
V[
p2496
tp2497
a(g423
Vline
p2498
tp2499
a(g693
g1417
tp2500
a(g826
g958
tp2501
a(g881
Vstring
p2502
tp2503
a(g693
g1417
tp2504
a(g826
g958
tp2505
a(g423
Vside
p2506
tp2507
a(g693
g1417
tp2508
a(g826
g958
tp2509
a(g423
Vwidth
p2510
tp2511
a(g693
V]
p2512
tp2513
a(g826
g958
tp2514
a(g693
g962
tp2515
a(g826
V\u000a
p2516
tp2517
a(g7
Vbegin
p2518
tp2519
a(g826
V\u000a
p2520
tp2521
a(g826
V    
p2522
tp2523
a(g423
Vswrite
p2524
tp2525
a(g693
g1018
tp2526
a(g423
Vmy_line
p2527
tp2528
a(g693
g1417
tp2529
a(g826
g958
tp2530
a(g76
V"sqrt( "
p2531
tp2532
a(g693
g1048
tp2533
a(g693
g962
tp2534
a(g826
V\u000a
p2535
tp2536
a(g826
V    
p2537
tp2538
a(g423
Vwrite
p2539
tp2540
a(g693
g1018
tp2541
a(g423
Vmy_line
p2542
tp2543
a(g693
g1417
tp2544
a(g826
g958
tp2545
a(g423
g2425
tp2546
a(g693
g1048
tp2547
a(g693
g962
tp2548
a(g826
V\u000a
p2549
tp2550
a(g826
V    
p2551
tp2552
a(g423
Vswrite
p2553
tp2554
a(g693
g1018
tp2555
a(g423
Vmy_line
p2556
tp2557
a(g693
g1417
tp2558
a(g826
g958
tp2559
a(g76
V" )= "
p2560
tp2561
a(g693
g1048
tp2562
a(g693
g962
tp2563
a(g826
V\u000a
p2564
tp2565
a(g826
V    
p2566
tp2567
a(g423
Vwrite
p2568
tp2569
a(g693
g1018
tp2570
a(g423
Vmy_line
p2571
tp2572
a(g693
g1417
tp2573
a(g826
g958
tp2574
a(g423
g2446
tp2575
a(g693
g1048
tp2576
a(g693
g962
tp2577
a(g826
V\u000a
p2578
tp2579
a(g826
V    
p2580
tp2581
a(g423
Vwriteline
p2582
tp2583
a(g693
g1018
tp2584
a(g423
Voutput
p2585
tp2586
a(g693
g1417
tp2587
a(g826
g958
tp2588
a(g423
Vmy_line
p2589
tp2590
a(g693
g1048
tp2591
a(g693
g962
tp2592
a(g826
V\u000a
p2593
tp2594
a(g7
Vend
p2595
tp2596
a(g826
g958
tp2597
a(g616
Vprint
p2598
tp2599
a(g693
g962
tp2600
a(g826
V\u000a
p2601
tp2602
a(g826
V\u000a
p2603
tp2604
a(g826
V\u000a
p2605
tp2606
a(g7
Ventity
p2607
tp2608
a(g826
g958
tp2609
a(g616
Vadd32csa
p2610
tp2611
a(g826
g958
tp2612
a(g7
Vis
p2613
tp2614
a(g826
V          
p2615
tp2616
a(g745
V-- one stage of carry save adder for multiplier
p2617
tp2618
a(g826
V\u000a
p2619
tp2620
a(g826
V  
p2621
tp2622
a(g7
Vport
p2623
tp2624
a(g693
g1018
tp2625
a(g826
V\u000a
p2626
tp2627
a(g826
V    
p2628
tp2629
a(g423
Vb
p2630
tp2631
a(g826
V       
p2632
tp2633
a(g400
g1030
tp2634
a(g826
g958
tp2635
a(g7
Vin
p2636
tp2637
a(g826
V  
p2638
tp2639
a(g881
Vstd_logic
p2640
tp2641
a(g693
g962
tp2642
a(g826
V                      
p2643
tp2644
a(g745
V-- a multiplier bit
p2645
tp2646
a(g826
V\u000a
p2647
tp2648
a(g826
V    
p2649
tp2650
a(g423
Va
p2651
tp2652
a(g826
V       
p2653
tp2654
a(g400
g1030
tp2655
a(g826
g958
tp2656
a(g7
Vin
p2657
tp2658
a(g826
V  
p2659
tp2660
a(g881
Vstd_logic_vector
p2661
tp2662
a(g693
g1018
tp2663
a(g22
V31
p2664
tp2665
a(g826
g958
tp2666
a(g7
Vdownto
p2667
tp2668
a(g826
g958
tp2669
a(g22
g1184
tp2670
a(g693
g1048
tp2671
a(g693
g962
tp2672
a(g826
V  
p2673
tp2674
a(g745
V-- multiplicand
p2675
tp2676
a(g826
V\u000a
p2677
tp2678
a(g826
V    
p2679
tp2680
a(g423
Vsum_in
p2681
tp2682
a(g826
V  
p2683
tp2684
a(g400
g1030
tp2685
a(g826
g958
tp2686
a(g7
Vin
p2687
tp2688
a(g826
V  
p2689
tp2690
a(g881
Vstd_logic_vector
p2691
tp2692
a(g693
g1018
tp2693
a(g22
V31
p2694
tp2695
a(g826
g958
tp2696
a(g7
Vdownto
p2697
tp2698
a(g826
g958
tp2699
a(g22
g1184
tp2700
a(g693
g1048
tp2701
a(g693
g962
tp2702
a(g826
V  
p2703
tp2704
a(g745
V-- sums from previous stage
p2705
tp2706
a(g826
V\u000a
p2707
tp2708
a(g826
V    
p2709
tp2710
a(g423
Vcin
p2711
tp2712
a(g826
V     
p2713
tp2714
a(g400
g1030
tp2715
a(g826
g958
tp2716
a(g7
Vin
p2717
tp2718
a(g826
V  
p2719
tp2720
a(g881
Vstd_logic_vector
p2721
tp2722
a(g693
g1018
tp2723
a(g22
V31
p2724
tp2725
a(g826
g958
tp2726
a(g7
Vdownto
p2727
tp2728
a(g826
g958
tp2729
a(g22
g1184
tp2730
a(g693
g1048
tp2731
a(g693
g962
tp2732
a(g826
V  
p2733
tp2734
a(g745
V-- carrys from previous stage
p2735
tp2736
a(g826
V\u000a
p2737
tp2738
a(g826
V    
p2739
tp2740
a(g423
Vsum_out
p2741
tp2742
a(g826
g958
tp2743
a(g400
g1030
tp2744
a(g826
g958
tp2745
a(g7
Vout
p2746
tp2747
a(g826
g958
tp2748
a(g881
Vstd_logic_vector
p2749
tp2750
a(g693
g1018
tp2751
a(g22
V31
p2752
tp2753
a(g826
g958
tp2754
a(g7
Vdownto
p2755
tp2756
a(g826
g958
tp2757
a(g22
g1184
tp2758
a(g693
g1048
tp2759
a(g693
g962
tp2760
a(g826
V  
p2761
tp2762
a(g745
V-- sums to next stage
p2763
tp2764
a(g826
V\u000a
p2765
tp2766
a(g826
V    
p2767
tp2768
a(g423
Vcout
p2769
tp2770
a(g826
V    
p2771
tp2772
a(g400
g1030
tp2773
a(g826
g958
tp2774
a(g7
Vout
p2775
tp2776
a(g826
g958
tp2777
a(g881
Vstd_logic_vector
p2778
tp2779
a(g693
g1018
tp2780
a(g22
V31
p2781
tp2782
a(g826
g958
tp2783
a(g7
Vdownto
p2784
tp2785
a(g826
g958
tp2786
a(g22
g1184
tp2787
a(g693
g1048
tp2788
a(g693
g1048
tp2789
a(g693
g962
tp2790
a(g826
g958
tp2791
a(g745
V-- carrys to next stage
p2792
tp2793
a(g826
V\u000a
p2794
tp2795
a(g7
Vend
p2796
tp2797
a(g826
g958
tp2798
a(g616
Vadd32csa
p2799
tp2800
a(g693
g962
tp2801
a(g826
V\u000a
p2802
tp2803
a(g826
V\u000a
p2804
tp2805
a(g826
V\u000a
p2806
tp2807
a(g7
VARCHITECTURE
p2808
tp2809
a(g826
g958
tp2810
a(g616
Vcircuits
p2811
tp2812
a(g826
g958
tp2813
a(g7
Vof
p2814
tp2815
a(g826
g958
tp2816
a(g616
Vadd32csa
p2817
tp2818
a(g826
g958
tp2819
a(g7
VIS
p2820
tp2821
a(g826
V\u000a
p2822
tp2823
a(g826
V  
p2824
tp2825
a(g7
VSIGNAL
p2826
tp2827
a(g826
g958
tp2828
a(g423
Vzero
p2829
tp2830
a(g826
g958
tp2831
a(g400
g1030
tp2832
a(g826
g958
tp2833
a(g881
VSTD_LOGIC_VECTOR
p2834
tp2835
a(g693
g1018
tp2836
a(g22
V31
p2837
tp2838
a(g826
g958
tp2839
a(g7
Vdownto
p2840
tp2841
a(g826
g958
tp2842
a(g22
g1184
tp2843
a(g693
g1048
tp2844
a(g826
g958
tp2845
a(g400
g1030
tp2846
a(g400
g1037
tp2847
a(g826
g958
tp2848
a(g285
VX"00000000"
p2849
tp2850
a(g693
g962
tp2851
a(g826
V\u000a
p2852
tp2853
a(g826
V  
p2854
tp2855
a(g7
VSIGNAL
p2856
tp2857
a(g826
g958
tp2858
a(g423
Vaa
p2859
tp2860
a(g826
g958
tp2861
a(g400
g1030
tp2862
a(g826
g958
tp2863
a(g881
Vstd_logic_vector
p2864
tp2865
a(g693
g1018
tp2866
a(g22
V31
p2867
tp2868
a(g826
g958
tp2869
a(g7
Vdownto
p2870
tp2871
a(g826
g958
tp2872
a(g22
g1184
tp2873
a(g693
g1048
tp2874
a(g826
g958
tp2875
a(g400
g1030
tp2876
a(g400
g1037
tp2877
a(g826
g958
tp2878
a(g285
VX"00000000"
p2879
tp2880
a(g693
g962
tp2881
a(g826
V\u000a
p2882
tp2883
a(g826
V  \u000a  
p2884
tp2885
a(g7
VCOMPONENT
p2886
tp2887
a(g826
g958
tp2888
a(g616
Vfadd
p2889
tp2890
a(g826
V    
p2891
tp2892
a(g745
V-- duplicates entity port
p2893
tp2894
a(g826
V\u000a
p2895
tp2896
a(g826
V    
p2897
tp2898
a(g7
VPoRT
p2899
tp2900
a(g693
g1018
tp2901
a(g423
g2651
tp2902
a(g826
V    
p2903
tp2904
a(g400
g1030
tp2905
a(g826
g958
tp2906
a(g7
Vin
p2907
tp2908
a(g826
V  
p2909
tp2910
a(g881
Vstd_logic
p2911
tp2912
a(g693
g962
tp2913
a(g826
V\u000a
p2914
tp2915
a(g826
V         
p2916
tp2917
a(g423
g2630
tp2918
a(g826
V    
p2919
tp2920
a(g400
g1030
tp2921
a(g826
g958
tp2922
a(g7
Vin
p2923
tp2924
a(g826
V  
p2925
tp2926
a(g881
Vstd_logic
p2927
tp2928
a(g693
g962
tp2929
a(g826
V\u000a
p2930
tp2931
a(g826
V         
p2932
tp2933
a(g423
Vcin
p2934
tp2935
a(g826
V  
p2936
tp2937
a(g400
g1030
tp2938
a(g826
g958
tp2939
a(g7
Vin
p2940
tp2941
a(g826
V  
p2942
tp2943
a(g881
Vstd_logic
p2944
tp2945
a(g693
g962
tp2946
a(g826
V\u000a
p2947
tp2948
a(g826
V         
p2949
tp2950
a(g423
Vs
p2951
tp2952
a(g826
V    
p2953
tp2954
a(g400
g1030
tp2955
a(g826
g958
tp2956
a(g7
Vout
p2957
tp2958
a(g826
g958
tp2959
a(g881
Vstd_logic
p2960
tp2961
a(g693
g962
tp2962
a(g826
V\u000a
p2963
tp2964
a(g826
V         
p2965
tp2966
a(g423
Vcout
p2967
tp2968
a(g826
g958
tp2969
a(g400
g1030
tp2970
a(g826
g958
tp2971
a(g7
Vout
p2972
tp2973
a(g826
g958
tp2974
a(g881
Vstd_logic
p2975
tp2976
a(g693
g1048
tp2977
a(g693
g962
tp2978
a(g826
V\u000a
p2979
tp2980
a(g826
V  
p2981
tp2982
a(g7
Vend
p2983
tp2984
a(g826
g958
tp2985
a(g7
VcomPonent
p2986
tp2987
a(g826
g958
tp2988
a(g616
Vfadd
p2989
tp2990
a(g693
g962
tp2991
a(g826
V\u000a
p2992
tp2993
a(g826
V  \u000a
p2994
tp2995
a(g7
Vbegin
p2996
tp2997
a(g826
V  
p2998
tp2999
a(g745
V-- circuits of add32csa
p3000
tp3001
a(g826
V\u000a
p3002
tp3003
a(g826
V  
p3004
tp3005
a(g423
Vaa
p3006
tp3007
a(g826
g958
tp3008
a(g400
g1630
tp3009
a(g400
g1037
tp3010
a(g826
g958
tp3011
a(g423
g2651
tp3012
a(g826
g958
tp3013
a(g7
Vwhen
p3014
tp3015
a(g826
g958
tp3016
a(g423
g2630
tp3017
a(g400
g1037
tp3018
a(g80
V'1'
p3019
tp3020
a(g826
g958
tp3021
a(g7
Velse
p3022
tp3023
a(g826
g958
tp3024
a(g423
Vzero
p3025
tp3026
a(g826
g958
tp3027
a(g7
Vafter
p3028
tp3029
a(g826
g958
tp3030
a(g22
g1178
tp3031
a(g826
g958
tp3032
a(g423
Vns
p3033
tp3034
a(g693
g962
tp3035
a(g826
V\u000a
p3036
tp3037
a(g826
V  
p3038
tp3039
a(g616
Vstage
p3040
tp3041
a(g400
g1030
tp3042
a(g826
g958
tp3043
a(g7
Vfor
p3044
tp3045
a(g826
g958
tp3046
a(g423
VI
p3047
tp3048
a(g826
g958
tp3049
a(g7
Vin
p3050
tp3051
a(g826
g958
tp3052
a(g22
g1184
tp3053
a(g826
g958
tp3054
a(g7
Vto
p3055
tp3056
a(g826
g958
tp3057
a(g22
V31
p3058
tp3059
a(g826
g958
tp3060
a(g7
Vgenerate
p3061
tp3062
a(g826
V\u000a
p3063
tp3064
a(g826
V    
p3065
tp3066
a(g423
Vsta
p3067
tp3068
a(g400
g1030
tp3069
a(g826
g958
tp3070
a(g423
Vfadd
p3071
tp3072
a(g826
g958
tp3073
a(g7
Vport
p3074
tp3075
a(g826
g958
tp3076
a(g7
Vmap
p3077
tp3078
a(g693
g1018
tp3079
a(g423
Vaa
p3080
tp3081
a(g693
g1018
tp3082
a(g423
g3047
tp3083
a(g693
g1048
tp3084
a(g693
g1417
tp3085
a(g826
g958
tp3086
a(g423
Vsum_in
p3087
tp3088
a(g693
g1018
tp3089
a(g423
g3047
tp3090
a(g693
g1048
tp3091
a(g693
g1417
tp3092
a(g826
g958
tp3093
a(g423
Vcin
p3094
tp3095
a(g693
g1018
tp3096
a(g423
g3047
tp3097
a(g693
g1048
tp3098
a(g826
g958
tp3099
a(g693
g1417
tp3100
a(g826
g958
tp3101
a(g423
Vsum_out
p3102
tp3103
a(g693
g1018
tp3104
a(g423
g3047
tp3105
a(g693
g1048
tp3106
a(g693
g1417
tp3107
a(g826
g958
tp3108
a(g423
Vcout
p3109
tp3110
a(g693
g1018
tp3111
a(g423
g3047
tp3112
a(g693
g1048
tp3113
a(g693
g1048
tp3114
a(g693
g962
tp3115
a(g826
V\u000a
p3116
tp3117
a(g826
V  
p3118
tp3119
a(g7
Vend
p3120
tp3121
a(g826
g958
tp3122
a(g7
Vgenerate
p3123
tp3124
a(g826
g958
tp3125
a(g616
Vstage
p3126
tp3127
a(g693
g962
tp3128
a(g826
V  \u000a
p3129
tp3130
a(g7
Vend
p3131
tp3132
a(g826
g958
tp3133
a(g7
Varchitecture
p3134
tp3135
a(g826
g958
tp3136
a(g616
Vcircuits
p3137
tp3138
a(g693
g962
tp3139
a(g826
g958
tp3140
a(g745
V-- of add32csa
p3141
tp3142
a(g826
V\u000a
p3143
tp3144
a.