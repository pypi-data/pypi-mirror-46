(lp0
(ccopy_reg
_reconstructor
p1
(cpygments.token
_TokenType
p2
c__builtin__
tuple
p3
(S'Comment'
p4
S'Preproc'
p5
tp6
tp7
Rp8
(dp9
S'parent'
p10
g1
(g2
g3
(g4
tp11
tp12
Rp13
(dp14
S'Multi'
p15
g1
(g2
g3
(g4
g15
tp16
tp17
Rp18
(dp19
g10
g13
sS'subtypes'
p20
c__builtin__
set
p21
((lp22
tp23
Rp24
sbsg10
g1
(g2
g3
(ttp25
Rp26
(dp27
S'Number'
p28
g1
(g2
g3
(S'Literal'
p29
g28
tp30
tp31
Rp32
(dp33
S'Integer'
p34
g1
(g2
g3
(g29
g28
g34
tp35
tp36
Rp37
(dp38
g10
g32
sS'Long'
p39
g1
(g2
g3
(g29
g28
g34
g39
tp40
tp41
Rp42
(dp43
g10
g37
sg20
g21
((lp44
tp45
Rp46
sbsg20
g21
((lp47
g42
atp48
Rp49
sbsg10
g1
(g2
g3
(g29
tp50
tp51
Rp52
(dp53
S'Scalar'
p54
g1
(g2
g3
(g29
g54
tp55
tp56
Rp57
(dp58
g10
g52
sg20
g21
((lp59
g1
(g2
g3
(g29
g54
S'Plain'
p60
tp61
tp62
Rp63
(dp64
g10
g57
sg20
g21
((lp65
tp66
Rp67
sbatp68
Rp69
sg60
g63
sbsg28
g32
sg10
g26
sS'Other'
p70
g1
(g2
g3
(g29
g70
tp71
tp72
Rp73
(dp74
g10
g52
sg20
g21
((lp75
tp76
Rp77
sbsS'Char'
p78
g1
(g2
g3
(g29
g78
tp79
tp80
Rp81
(dp82
g10
g52
sg20
g21
((lp83
tp84
Rp85
sbsS'String'
p86
g1
(g2
g3
(g29
g86
tp87
tp88
Rp89
(dp90
g78
g1
(g2
g3
(g29
g86
g78
tp91
tp92
Rp93
(dp94
g10
g89
sg20
g21
((lp95
tp96
Rp97
sbsS'Backtick'
p98
g1
(g2
g3
(g29
g86
g98
tp99
tp100
Rp101
(dp102
g10
g89
sg20
g21
((lp103
tp104
Rp105
sbsS'Heredoc'
p106
g1
(g2
g3
(g29
g86
g106
tp107
tp108
Rp109
(dp110
g10
g89
sg20
g21
((lp111
tp112
Rp113
sbsS'Symbol'
p114
g1
(g2
g3
(g29
g86
g114
tp115
tp116
Rp117
(dp118
g10
g89
sg20
g21
((lp119
tp120
Rp121
sbsS'Interpol'
p122
g1
(g2
g3
(g29
g86
g122
tp123
tp124
Rp125
(dp126
g10
g89
sg20
g21
((lp127
tp128
Rp129
sbsS'Delimiter'
p130
g1
(g2
g3
(g29
g86
g130
tp131
tp132
Rp133
(dp134
g10
g89
sg20
g21
((lp135
tp136
Rp137
sbsS'Boolean'
p138
g1
(g2
g3
(g29
g86
g138
tp139
tp140
Rp141
(dp142
g10
g89
sg20
g21
((lp143
tp144
Rp145
sbsS'Character'
p146
g1
(g2
g3
(g29
g86
g146
tp147
tp148
Rp149
(dp150
g10
g89
sg20
g21
((lp151
tp152
Rp153
sbsS'Double'
p154
g1
(g2
g3
(g29
g86
g154
tp155
tp156
Rp157
(dp158
g10
g89
sg20
g21
((lp159
tp160
Rp161
sbsS'Delimeter'
p162
g1
(g2
g3
(g29
g86
g162
tp163
tp164
Rp165
(dp166
g10
g89
sg20
g21
((lp167
tp168
Rp169
sbsS'Atom'
p170
g1
(g2
g3
(g29
g86
g170
tp171
tp172
Rp173
(dp174
g10
g89
sg20
g21
((lp175
tp176
Rp177
sbsS'Affix'
p178
g1
(g2
g3
(g29
g86
g178
tp179
tp180
Rp181
(dp182
g10
g89
sg20
g21
((lp183
tp184
Rp185
sbsS'Name'
p186
g1
(g2
g3
(g29
g86
g186
tp187
tp188
Rp189
(dp190
g10
g89
sg20
g21
((lp191
tp192
Rp193
sbsS'Regex'
p194
g1
(g2
g3
(g29
g86
g194
tp195
tp196
Rp197
(dp198
g10
g89
sg20
g21
((lp199
tp200
Rp201
sbsS'Interp'
p202
g1
(g2
g3
(g29
g86
g202
tp203
tp204
Rp205
(dp206
g10
g89
sg20
g21
((lp207
tp208
Rp209
sbsS'Escape'
p210
g1
(g2
g3
(g29
g86
g210
tp211
tp212
Rp213
(dp214
g10
g89
sg20
g21
((lp215
tp216
Rp217
sbsg20
g21
((lp218
g133
ag117
ag197
ag1
(g2
g3
(g29
g86
S'Doc'
p219
tp220
tp221
Rp222
(dp223
g10
g89
sg20
g21
((lp224
tp225
Rp226
sbag149
ag141
ag157
ag125
ag173
ag165
ag189
ag213
ag1
(g2
g3
(g29
g86
S'Single'
p227
tp228
tp229
Rp230
(dp231
g10
g89
sg20
g21
((lp232
tp233
Rp234
sbag1
(g2
g3
(g29
g86
g70
tp235
tp236
Rp237
(dp238
g10
g89
sg20
g21
((lp239
tp240
Rp241
sbag205
ag101
ag181
ag1
(g2
g3
(g29
g86
S'Moment'
p242
tp243
tp244
Rp245
(dp246
g10
g89
sg20
g21
((lp247
tp248
Rp249
sbag93
ag109
atp250
Rp251
sg227
g230
sg242
g245
sg10
g52
sg70
g237
sg219
g222
sbsg20
g21
((lp252
g89
ag81
ag73
ag1
(g2
g3
(g29
S'Date'
p253
tp254
tp255
Rp256
(dp257
g10
g52
sg20
g21
((lp258
tp259
Rp260
sbag57
ag32
atp261
Rp262
sg253
g256
sbsS'Bin'
p263
g1
(g2
g3
(g29
g28
g263
tp264
tp265
Rp266
(dp267
g10
g32
sg20
g21
((lp268
tp269
Rp270
sbsS'Radix'
p271
g1
(g2
g3
(g29
g28
g271
tp272
tp273
Rp274
(dp275
g10
g32
sg20
g21
((lp276
tp277
Rp278
sbsS'Oct'
p279
g1
(g2
g3
(g29
g28
g279
tp280
tp281
Rp282
(dp283
g10
g32
sg20
g21
((lp284
tp285
Rp286
sbsS'Dec'
p287
g1
(g2
g3
(g29
g28
g287
tp288
tp289
Rp290
(dp291
g10
g32
sg20
g21
((lp292
tp293
Rp294
sbsS'Hex'
p295
g1
(g2
g3
(g29
g28
g295
tp296
tp297
Rp298
(dp299
g10
g32
sg20
g21
((lp300
tp301
Rp302
sbsg20
g21
((lp303
g37
ag274
ag290
ag1
(g2
g3
(g29
g28
S'Decimal'
p304
tp305
tp306
Rp307
(dp308
g10
g32
sg20
g21
((lp309
tp310
Rp311
sbag266
ag1
(g2
g3
(g29
g28
S'Float'
p312
tp313
tp314
Rp315
(dp316
g10
g32
sg20
g21
((lp317
tp318
Rp319
sbag282
ag298
atp320
Rp321
sg304
g307
sg312
g315
sbsS'Generic'
p322
g1
(g2
g3
(g322
tp323
tp324
Rp325
(dp326
g10
g26
sS'Deleted'
p327
g1
(g2
g3
(g322
g327
tp328
tp329
Rp330
(dp331
g10
g325
sg20
g21
((lp332
tp333
Rp334
sbsS'Subheading'
p335
g1
(g2
g3
(g322
g335
tp336
tp337
Rp338
(dp339
g10
g325
sg20
g21
((lp340
tp341
Rp342
sbsS'Heading'
p343
g1
(g2
g3
(g322
g343
tp344
tp345
Rp346
(dp347
g10
g325
sg20
g21
((lp348
tp349
Rp350
sbsS'Emph'
p351
g1
(g2
g3
(g322
g351
tp352
tp353
Rp354
(dp355
g10
g325
sg20
g21
((lp356
tp357
Rp358
sbsS'Prompt'
p359
g1
(g2
g3
(g322
g359
tp360
tp361
Rp362
(dp363
g10
g325
sg20
g21
((lp364
tp365
Rp366
sbsS'Inserted'
p367
g1
(g2
g3
(g322
g367
tp368
tp369
Rp370
(dp371
g10
g325
sg20
g21
((lp372
tp373
Rp374
sbsS'Strong'
p375
g1
(g2
g3
(g322
g375
tp376
tp377
Rp378
(dp379
g10
g325
sg20
g21
((lp380
tp381
Rp382
sbsS'Error'
p383
g1
(g2
g3
(g322
g383
tp384
tp385
Rp386
(dp387
g10
g325
sg20
g21
((lp388
tp389
Rp390
sbsS'Traceback'
p391
g1
(g2
g3
(g322
g391
tp392
tp393
Rp394
(dp395
g10
g325
sg20
g21
((lp396
tp397
Rp398
sbsg20
g21
((lp399
g346
ag338
ag1
(g2
g3
(g322
S'Output'
p400
tp401
tp402
Rp403
(dp404
g10
g325
sg20
g21
((lp405
tp406
Rp407
sbag378
ag354
ag386
ag394
ag370
ag362
ag330
atp408
Rp409
sg400
g403
sbsS'Operator'
p410
g1
(g2
g3
(g410
tp411
tp412
Rp413
(dp414
g10
g26
sS'DBS'
p415
g1
(g2
g3
(g410
g415
tp416
tp417
Rp418
(dp419
g10
g413
sg20
g21
((lp420
tp421
Rp422
sbsg20
g21
((lp423
g418
ag1
(g2
g3
(g410
S'Word'
p424
tp425
tp426
Rp427
(dp428
g10
g413
sg20
g21
((lp429
tp430
Rp431
sbatp432
Rp433
sg424
g427
sbsg86
g89
sg186
g1
(g2
g3
(g186
tp434
tp435
Rp436
(dp437
S'Variable'
p438
g1
(g2
g3
(g186
g438
tp439
tp440
Rp441
(dp442
g10
g436
sS'Class'
p443
g1
(g2
g3
(g186
g438
g443
tp444
tp445
Rp446
(dp447
g10
g441
sg20
g21
((lp448
tp449
Rp450
sbsS'Anonymous'
p451
g1
(g2
g3
(g186
g438
g451
tp452
tp453
Rp454
(dp455
g10
g441
sg20
g21
((lp456
tp457
Rp458
sbsS'Instance'
p459
g1
(g2
g3
(g186
g438
g459
tp460
tp461
Rp462
(dp463
g10
g441
sg20
g21
((lp464
tp465
Rp466
sbsS'Global'
p467
g1
(g2
g3
(g186
g438
g467
tp468
tp469
Rp470
(dp471
g10
g441
sg20
g21
((lp472
tp473
Rp474
sbsg20
g21
((lp475
g454
ag462
ag1
(g2
g3
(g186
g438
S'Magic'
p476
tp477
tp478
Rp479
(dp480
g10
g441
sg20
g21
((lp481
tp482
Rp483
sbag470
ag446
atp484
Rp485
sg476
g479
sbsg410
g1
(g2
g3
(g186
g410
tp486
tp487
Rp488
(dp489
g10
g436
sg20
g21
((lp490
tp491
Rp492
sbsS'Decorator'
p493
g1
(g2
g3
(g186
g493
tp494
tp495
Rp496
(dp497
g10
g436
sg20
g21
((lp498
tp499
Rp500
sbsS'Entity'
p501
g1
(g2
g3
(g186
g501
tp502
tp503
Rp504
(dp505
g10
g436
sg415
g1
(g2
g3
(g186
g501
g415
tp506
tp507
Rp508
(dp509
g10
g504
sg20
g21
((lp510
tp511
Rp512
sbsg20
g21
((lp513
g508
atp514
Rp515
sbsg114
g1
(g2
g3
(g186
g114
tp516
tp517
Rp518
(dp519
g10
g436
sg20
g21
((lp520
tp521
Rp522
sbsS'Property'
p523
g1
(g2
g3
(g186
g523
tp524
tp525
Rp526
(dp527
g10
g436
sg20
g21
((lp528
tp529
Rp530
sbsS'Pseudo'
p531
g1
(g2
g3
(g186
g531
tp532
tp533
Rp534
(dp535
g10
g436
sg20
g21
((lp536
tp537
Rp538
sbsS'Type'
p539
g1
(g2
g3
(g186
g539
tp540
tp541
Rp542
(dp543
g10
g436
sg20
g21
((lp544
tp545
Rp546
sbsS'Classes'
p547
g1
(g2
g3
(g186
g547
tp548
tp549
Rp550
(dp551
g10
g436
sg20
g21
((lp552
tp553
Rp554
sbsS'Tag'
p555
g1
(g2
g3
(g186
g555
tp556
tp557
Rp558
(dp559
g10
g436
sg20
g21
((lp560
tp561
Rp562
sbsS'Constant'
p563
g1
(g2
g3
(g186
g563
tp564
tp565
Rp566
(dp567
g10
g436
sg20
g21
((lp568
tp569
Rp570
sbsS'Function'
p571
g1
(g2
g3
(g186
g571
tp572
tp573
Rp574
(dp575
g10
g436
sg20
g21
((lp576
g1
(g2
g3
(g186
g571
g476
tp577
tp578
Rp579
(dp580
g10
g574
sg20
g21
((lp581
tp582
Rp583
sbatp584
Rp585
sg476
g579
sbsS'Blubb'
p586
g1
(g2
g3
(g186
g586
tp587
tp588
Rp589
(dp590
g10
g436
sg20
g21
((lp591
tp592
Rp593
sbsS'Label'
p594
g1
(g2
g3
(g186
g594
tp595
tp596
Rp597
(dp598
g10
g436
sg20
g21
((lp599
tp600
Rp601
sbsS'Field'
p602
g1
(g2
g3
(g186
g602
tp603
tp604
Rp605
(dp606
g10
g436
sg20
g21
((lp607
tp608
Rp609
sbsS'Exception'
p610
g1
(g2
g3
(g186
g610
tp611
tp612
Rp613
(dp614
g10
g436
sg20
g21
((lp615
tp616
Rp617
sbsS'Namespace'
p618
g1
(g2
g3
(g186
g618
tp619
tp620
Rp621
(dp622
g10
g436
sg20
g21
((lp623
tp624
Rp625
sbsg20
g21
((lp626
g496
ag589
ag534
ag504
ag441
ag613
ag526
ag558
ag574
ag550
ag1
(g2
g3
(g186
g443
tp627
tp628
Rp629
(dp630
g10
g436
sg415
g1
(g2
g3
(g186
g443
g415
tp631
tp632
Rp633
(dp634
g10
g629
sg20
g21
((lp635
tp636
Rp637
sbsg20
g21
((lp638
g1
(g2
g3
(g186
g443
S'Start'
p639
tp640
tp641
Rp642
(dp643
g10
g629
sg20
g21
((lp644
tp645
Rp646
sbag633
atp647
Rp648
sg639
g642
sbag1
(g2
g3
(g186
g70
tp649
tp650
Rp651
(dp652
g10
g436
sS'Member'
p653
g1
(g2
g3
(g186
g70
g653
tp654
tp655
Rp656
(dp657
g10
g651
sg20
g21
((lp658
tp659
Rp660
sbsg20
g21
((lp661
g656
atp662
Rp663
sbag597
ag488
ag621
ag1
(g2
g3
(g186
S'Attribute'
p664
tp665
tp666
Rp667
(dp668
g10
g436
sg438
g1
(g2
g3
(g186
g664
g438
tp669
tp670
Rp671
(dp672
g10
g667
sg20
g21
((lp673
tp674
Rp675
sbsg20
g21
((lp676
g671
atp677
Rp678
sbag566
ag1
(g2
g3
(g186
S'Builtin'
p679
tp680
tp681
Rp682
(dp683
g10
g436
sg539
g1
(g2
g3
(g186
g679
g539
tp684
tp685
Rp686
(dp687
g10
g682
sg20
g21
((lp688
tp689
Rp690
sbsg20
g21
((lp691
g1
(g2
g3
(g186
g679
g531
tp692
tp693
Rp694
(dp695
g10
g682
sg20
g21
((lp696
tp697
Rp698
sbag686
atp699
Rp700
sg531
g694
sbag605
ag542
ag518
atp701
Rp702
sg10
g26
sg443
g629
sg679
g682
sg664
g667
sg70
g651
sbsS'Punctuation'
p703
g1
(g2
g3
(g703
tp704
tp705
Rp706
(dp707
g10
g26
sg20
g21
((lp708
g1
(g2
g3
(g703
S'Indicator'
p709
tp710
tp711
Rp712
(dp713
g10
g706
sg20
g21
((lp714
tp715
Rp716
sbatp717
Rp718
sg709
g712
sbsg4
g13
sg29
g52
sg70
g1
(g2
g3
(g70
tp719
tp720
Rp721
(dp722
g10
g26
sg20
g21
((lp723
tp724
Rp725
sbsg383
g1
(g2
g3
(g383
tp726
tp727
Rp728
(dp729
g10
g26
sg20
g21
((lp730
tp731
Rp732
sbsS'Token'
p733
g26
sg210
g1
(g2
g3
(g210
tp734
tp735
Rp736
(dp737
g10
g26
sg20
g21
((lp738
tp739
Rp740
sbsg20
g21
((lp741
g436
ag721
ag1
(g2
g3
(S'Keyword'
p742
tp743
tp744
Rp745
(dp746
g10
g26
sg539
g1
(g2
g3
(g742
g539
tp747
tp748
Rp749
(dp750
g10
g745
sg20
g21
((lp751
tp752
Rp753
sbsS'Control'
p754
g1
(g2
g3
(g742
g754
tp755
tp756
Rp757
(dp758
g10
g745
sg20
g21
((lp759
tp760
Rp761
sbsg563
g1
(g2
g3
(g742
g563
tp762
tp763
Rp764
(dp765
g10
g745
sg20
g21
((lp766
tp767
Rp768
sbsg618
g1
(g2
g3
(g742
g618
tp769
tp770
Rp771
(dp772
g10
g745
sg20
g21
((lp773
tp774
Rp775
sbsS'PreProc'
p776
g1
(g2
g3
(g742
g776
tp777
tp778
Rp779
(dp780
g10
g745
sg20
g21
((lp781
tp782
Rp783
sbsg531
g1
(g2
g3
(g742
g531
tp784
tp785
Rp786
(dp787
g10
g745
sg20
g21
((lp788
tp789
Rp790
sbsS'Reserved'
p791
g1
(g2
g3
(g742
g791
tp792
tp793
Rp794
(dp795
g10
g745
sg20
g21
((lp796
tp797
Rp798
sbsg20
g21
((lp799
g771
ag1
(g2
g3
(g742
g424
tp800
tp801
Rp802
(dp803
g10
g745
sg20
g21
((lp804
tp805
Rp806
sbag757
ag1
(g2
g3
(g742
S'Declaration'
p807
tp808
tp809
Rp810
(dp811
g10
g745
sg20
g21
((lp812
tp813
Rp814
sbag1
(g2
g3
(g742
g742
tp815
tp816
Rp817
(dp818
g10
g745
sg20
g21
((lp819
tp820
Rp821
sbag786
ag764
ag749
ag794
ag779
atp822
Rp823
sg742
g817
sg807
g810
sg424
g802
sbag325
ag1
(g2
g3
(S'Text'
p824
tp825
tp826
Rp827
(dp828
S'Beer'
p829
g1
(g2
g3
(g824
g829
tp830
tp831
Rp832
(dp833
g10
g827
sg20
g21
((lp834
tp835
Rp836
sbsS'Whitespace'
p837
g1
(g2
g3
(g824
g837
tp838
tp839
Rp840
(dp841
g10
g827
sg20
g21
((lp842
tp843
Rp844
sbsg10
g26
sS'Root'
p845
g1
(g2
g3
(g824
g845
tp846
tp847
Rp848
(dp849
g10
g827
sg20
g21
((lp850
tp851
Rp852
sbsg114
g1
(g2
g3
(g824
g114
tp853
tp854
Rp855
(dp856
g10
g827
sg20
g21
((lp857
tp858
Rp859
sbsg703
g1
(g2
g3
(g824
g703
tp860
tp861
Rp862
(dp863
g10
g827
sg20
g21
((lp864
tp865
Rp866
sbsg20
g21
((lp867
g848
ag855
ag862
ag840
ag832
ag1
(g2
g3
(g824
S'Rag'
p868
tp869
tp870
Rp871
(dp872
g10
g827
sg20
g21
((lp873
tp874
Rp875
sbatp876
Rp877
sg868
g871
sbag413
ag736
ag706
ag13
ag728
ag52
atp878
Rp879
sg742
g745
sg824
g827
sbsS'Special'
p880
g1
(g2
g3
(g4
g880
tp881
tp882
Rp883
(dp884
g10
g13
sg20
g21
((lp885
tp886
Rp887
sbsS'Hashbang'
p888
g1
(g2
g3
(g4
g888
tp889
tp890
Rp891
(dp892
g10
g13
sg20
g21
((lp893
tp894
Rp895
sbsg5
g8
sg227
g1
(g2
g3
(g4
g227
tp896
tp897
Rp898
(dp899
g10
g13
sg20
g21
((lp900
tp901
Rp902
sbsS'Directive'
p903
g1
(g2
g3
(g4
g903
tp904
tp905
Rp906
(dp907
g10
g13
sg20
g21
((lp908
tp909
Rp910
sbsg219
g1
(g2
g3
(g4
g219
tp911
tp912
Rp913
(dp914
g10
g13
sg20
g21
((lp915
tp916
Rp917
sbsS'Singleline'
p918
g1
(g2
g3
(g4
g918
tp919
tp920
Rp921
(dp922
g10
g13
sg20
g21
((lp923
tp924
Rp925
sbsS'Multiline'
p926
g1
(g2
g3
(g4
g926
tp927
tp928
Rp929
(dp930
g10
g13
sg20
g21
((lp931
tp932
Rp933
sbsg20
g21
((lp934
g913
ag906
ag891
ag18
ag921
ag8
ag929
ag898
ag1
(g2
g3
(g4
S'PreprocFile'
p935
tp936
tp937
Rp938
(dp939
g10
g13
sg20
g21
((lp940
tp941
Rp942
sbag1
(g2
g3
(g4
S'SingleLine'
p943
tp944
tp945
Rp946
(dp947
g10
g13
sg20
g21
((lp948
tp949
Rp950
sbag883
atp951
Rp952
sg935
g938
sg943
g946
sbsg20
g21
((lp953
tp954
Rp955
sbV#ifdef ARCH_ARM\u000a
p956
tp957
a(g745
Varch
p958
tp959
a(g827
V 
p960
tp961
a(g745
Varm11
p962
tp963
a(g827
V\u000a
p964
tp965
a(g8
V#else\u000a
p966
tp967
a(g745
Varch
p968
tp969
a(g827
g960
tp970
a(g745
Via32
p971
tp972
a(g827
V\u000a
p973
tp974
a(g8
V#endif\u000a
p975
tp976
a(g827
V\u000a
p977
tp978
a(g745
Vobjects
p979
tp980
a(g827
g960
tp981
a(g706
V{
p982
tp983
a(g827
V\u000a  
p984
tp985
a(g436
Vmy_ep
p986
tp987
a(g827
g960
tp988
a(g706
V=
p989
tp990
a(g827
g960
tp991
a(g749
Vep
p992
tp993
a(g827
g960
tp994
a(g13
V/* A synchronous endpoint */
p995
tp996
a(g827
V\u000a\u000a  
p997
tp998
a(g13
V/* Two thread control blocks */
p999
tp1000
a(g827
V\u000a  
p1001
tp1002
a(g436
Vtcb1
p1003
tp1004
a(g827
g960
tp1005
a(g706
g989
tp1006
a(g827
g960
tp1007
a(g749
Vtcb
p1008
tp1009
a(g827
V\u000a  
p1010
tp1011
a(g436
Vtcb2
p1012
tp1013
a(g827
g960
tp1014
a(g706
g989
tp1015
a(g827
g960
tp1016
a(g749
Vtcb
p1017
tp1018
a(g827
V\u000a\u000a  
p1019
tp1020
a(g13
V/* Four frames of physical memory */
p1021
tp1022
a(g827
V\u000a  
p1023
tp1024
a(g436
Vframe1
p1025
tp1026
a(g827
g960
tp1027
a(g706
g989
tp1028
a(g827
g960
tp1029
a(g749
Vframe
p1030
tp1031
a(g827
g960
tp1032
a(g706
V(
p1033
tp1034
a(g32
V4k
p1035
tp1036
a(g706
V)
p1037
tp1038
a(g827
V\u000a  
p1039
tp1040
a(g436
Vframe2
p1041
tp1042
a(g827
g960
tp1043
a(g706
g989
tp1044
a(g827
g960
tp1045
a(g749
Vframe
p1046
tp1047
a(g827
g960
tp1048
a(g706
g1033
tp1049
a(g32
V4k
p1050
tp1051
a(g706
g1037
tp1052
a(g827
V\u000a  
p1053
tp1054
a(g436
Vframe3
p1055
tp1056
a(g827
g960
tp1057
a(g706
g989
tp1058
a(g827
g960
tp1059
a(g749
Vframe
p1060
tp1061
a(g827
g960
tp1062
a(g706
g1033
tp1063
a(g32
V4k
p1064
tp1065
a(g706
g1037
tp1066
a(g827
V\u000a  
p1067
tp1068
a(g436
Vframe4
p1069
tp1070
a(g827
g960
tp1071
a(g706
g989
tp1072
a(g827
g960
tp1073
a(g749
Vframe
p1074
tp1075
a(g827
g960
tp1076
a(g706
g1033
tp1077
a(g32
V4k
p1078
tp1079
a(g706
g1037
tp1080
a(g827
V\u000a\u000a  
p1081
tp1082
a(g13
V/* Two page tables */
p1083
tp1084
a(g827
V\u000a  
p1085
tp1086
a(g436
Vpt1
p1087
tp1088
a(g827
g960
tp1089
a(g706
g989
tp1090
a(g827
g960
tp1091
a(g749
Vpt
p1092
tp1093
a(g827
V\u000a  
p1094
tp1095
a(g436
Vpt2
p1096
tp1097
a(g827
g960
tp1098
a(g706
g989
tp1099
a(g827
g960
tp1100
a(g749
Vpt
p1101
tp1102
a(g827
V\u000a\u000a  
p1103
tp1104
a(g13
V/* Two page directories */
p1105
tp1106
a(g827
V\u000a  
p1107
tp1108
a(g436
Vpd1
p1109
tp1110
a(g827
g960
tp1111
a(g706
g989
tp1112
a(g827
g960
tp1113
a(g749
Vpd
p1114
tp1115
a(g827
V\u000a  
p1116
tp1117
a(g436
Vpd2
p1118
tp1119
a(g827
g960
tp1120
a(g706
g989
tp1121
a(g827
g960
tp1122
a(g749
Vpd
p1123
tp1124
a(g827
V\u000a\u000a  
p1125
tp1126
a(g13
V/* Two capability nodes */
p1127
tp1128
a(g827
V\u000a  
p1129
tp1130
a(g436
Vcnode1
p1131
tp1132
a(g827
g960
tp1133
a(g706
g989
tp1134
a(g827
g960
tp1135
a(g749
Vcnode
p1136
tp1137
a(g827
g960
tp1138
a(g706
g1033
tp1139
a(g32
V2
p1140
tp1141
a(g827
g960
tp1142
a(g32
Vbits
p1143
tp1144
a(g706
g1037
tp1145
a(g827
V\u000a  
p1146
tp1147
a(g436
Vcnode2
p1148
tp1149
a(g827
g960
tp1150
a(g706
g989
tp1151
a(g827
g960
tp1152
a(g749
Vcnode
p1153
tp1154
a(g827
g960
tp1155
a(g706
g1033
tp1156
a(g32
V3
p1157
tp1158
a(g827
g960
tp1159
a(g32
Vbits
p1160
tp1161
a(g706
g1037
tp1162
a(g827
V\u000a
p1163
tp1164
a(g706
V}
p1165
tp1166
a(g827
V\u000a
p1167
tp1168
a(g745
Vcaps
p1169
tp1170
a(g827
g960
tp1171
a(g706
g982
tp1172
a(g827
V\u000a  
p1173
tp1174
a(g436
Vcnode1
p1175
tp1176
a(g827
g960
tp1177
a(g706
g982
tp1178
a(g827
V\u000a    
p1179
tp1180
a(g298
V0x1
p1181
tp1182
a(g706
V:
p1183
tp1184
a(g827
g960
tp1185
a(g436
Vframe1
p1186
tp1187
a(g827
g960
tp1188
a(g706
g1033
tp1189
a(g794
VRW
p1190
tp1191
a(g706
g1037
tp1192
a(g827
g960
tp1193
a(g13
V/* read/write */
p1194
tp1195
a(g827
V\u000a    
p1196
tp1197
a(g298
V0x2
p1198
tp1199
a(g706
g1183
tp1200
a(g827
g960
tp1201
a(g436
Vmy_ep
p1202
tp1203
a(g827
g960
tp1204
a(g706
g1033
tp1205
a(g794
VR
p1206
tp1207
a(g706
g1037
tp1208
a(g827
V   
p1209
tp1210
a(g13
V/* read-only */
p1211
tp1212
a(g827
V\u000a  
p1213
tp1214
a(g706
g1165
tp1215
a(g827
V\u000a  
p1216
tp1217
a(g436
Vcnode2
p1218
tp1219
a(g827
g960
tp1220
a(g706
g982
tp1221
a(g827
V\u000a    
p1222
tp1223
a(g298
V0x1
p1224
tp1225
a(g706
g1183
tp1226
a(g827
g960
tp1227
a(g436
Vmy_ep
p1228
tp1229
a(g827
g960
tp1230
a(g706
g1033
tp1231
a(g794
VW
p1232
tp1233
a(g706
g1037
tp1234
a(g827
V   
p1235
tp1236
a(g13
V/* write-only */
p1237
tp1238
a(g827
V\u000a  
p1239
tp1240
a(g706
g1165
tp1241
a(g827
V\u000a  
p1242
tp1243
a(g436
Vtcb1
p1244
tp1245
a(g827
g960
tp1246
a(g706
g982
tp1247
a(g827
V\u000a    
p1248
tp1249
a(g32
Vvspace
p1250
tp1251
a(g706
g1183
tp1252
a(g827
g960
tp1253
a(g436
Vpd1
p1254
tp1255
a(g827
V\u000a    
p1256
tp1257
a(g32
Vipc_buffer_slot
p1258
tp1259
a(g706
g1183
tp1260
a(g827
g960
tp1261
a(g436
Vframe1
p1262
tp1263
a(g827
V\u000a    
p1264
tp1265
a(g32
Vcspace
p1266
tp1267
a(g706
g1183
tp1268
a(g827
g960
tp1269
a(g436
Vcnode1
p1270
tp1271
a(g827
V\u000a  
p1272
tp1273
a(g706
g1165
tp1274
a(g827
V\u000a  
p1275
tp1276
a(g436
Vpd1
p1277
tp1278
a(g827
g960
tp1279
a(g706
g982
tp1280
a(g827
V\u000a    
p1281
tp1282
a(g298
V0x10
p1283
tp1284
a(g706
g1183
tp1285
a(g827
g960
tp1286
a(g436
Vpt1
p1287
tp1288
a(g827
V\u000a  
p1289
tp1290
a(g706
g1165
tp1291
a(g827
V\u000a  
p1292
tp1293
a(g436
Vpt1
p1294
tp1295
a(g827
g960
tp1296
a(g706
g982
tp1297
a(g827
V\u000a    
p1298
tp1299
a(g298
V0x8
p1300
tp1301
a(g706
g1183
tp1302
a(g827
g960
tp1303
a(g436
Vframe1
p1304
tp1305
a(g827
g960
tp1306
a(g706
g1033
tp1307
a(g794
VRW
p1308
tp1309
a(g706
g1037
tp1310
a(g827
V\u000a    
p1311
tp1312
a(g298
V0x9
p1313
tp1314
a(g706
g1183
tp1315
a(g827
g960
tp1316
a(g436
Vframe2
p1317
tp1318
a(g827
g960
tp1319
a(g706
g1033
tp1320
a(g794
g1206
tp1321
a(g706
g1037
tp1322
a(g827
V\u000a  
p1323
tp1324
a(g706
g1165
tp1325
a(g827
V\u000a  
p1326
tp1327
a(g436
Vtcb2
p1328
tp1329
a(g827
g960
tp1330
a(g706
g982
tp1331
a(g827
V\u000a    
p1332
tp1333
a(g32
Vvspace
p1334
tp1335
a(g706
g1183
tp1336
a(g827
g960
tp1337
a(g436
Vpd2
p1338
tp1339
a(g827
V\u000a    
p1340
tp1341
a(g32
Vipc_buffer_slot
p1342
tp1343
a(g706
g1183
tp1344
a(g827
g960
tp1345
a(g436
Vframe3
p1346
tp1347
a(g827
V\u000a    
p1348
tp1349
a(g32
Vcspace
p1350
tp1351
a(g706
g1183
tp1352
a(g827
g960
tp1353
a(g436
Vcnode2
p1354
tp1355
a(g827
V\u000a  
p1356
tp1357
a(g706
g1165
tp1358
a(g827
V\u000a  
p1359
tp1360
a(g436
Vpd2
p1361
tp1362
a(g827
g960
tp1363
a(g706
g982
tp1364
a(g827
V\u000a    
p1365
tp1366
a(g298
V0x10
p1367
tp1368
a(g706
g1183
tp1369
a(g827
g960
tp1370
a(g436
Vpt2
p1371
tp1372
a(g827
V\u000a  
p1373
tp1374
a(g706
g1165
tp1375
a(g827
V\u000a  
p1376
tp1377
a(g436
Vpt2
p1378
tp1379
a(g827
g960
tp1380
a(g706
g982
tp1381
a(g827
V\u000a    
p1382
tp1383
a(g298
V0x10
p1384
tp1385
a(g706
g1183
tp1386
a(g827
g960
tp1387
a(g436
Vframe3
p1388
tp1389
a(g827
g960
tp1390
a(g706
g1033
tp1391
a(g794
VRW
p1392
tp1393
a(g706
g1037
tp1394
a(g827
V\u000a    
p1395
tp1396
a(g298
V0x12
p1397
tp1398
a(g706
g1183
tp1399
a(g827
g960
tp1400
a(g436
Vframe4
p1401
tp1402
a(g827
g960
tp1403
a(g706
g1033
tp1404
a(g794
g1206
tp1405
a(g706
g1037
tp1406
a(g827
V\u000a  
p1407
tp1408
a(g706
g1165
tp1409
a(g827
V\u000a
p1410
tp1411
a(g706
g1165
tp1412
a(g827
V\u000a
p1413
tp1414
a.